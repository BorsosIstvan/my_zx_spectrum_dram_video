//Copyright (C)2014-2025 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.11.03 Education
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9
//Device Version: C
//Created Time: Sun Sep 14 09:39:08 2025

module Gowin_pROM_0 (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [12:0] ad;

wire [29:0] prom_inst_0_dout_w;
wire [29:0] prom_inst_1_dout_w;
wire [29:0] prom_inst_2_dout_w;
wire [29:0] prom_inst_3_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[29:0],dout[1:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 2;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h1986C65551025FFFE71D165D56D507102C25AD19FFFFFF010586FFDBC3867FDF;
defparam prom_inst_0.INIT_RAM_01 = 256'h98E2323B67539BE7241887DB64FE79064F069060496F272905E4AD1BD2B32086;
defparam prom_inst_0.INIT_RAM_02 = 256'hCD02601E6DE690DA34A44E539C59999E5C7CF24DD96D16E1E8904F241921909B;
defparam prom_inst_0.INIT_RAM_03 = 256'h91A53D8CE597266798C0987C067504341C12673F0FB965164BE4BB66CD91058C;
defparam prom_inst_0.INIT_RAM_04 = 256'hDB3B274B07ADE12CF6D49F9EB1F221765A6B13D0035412F9C81C77A36AC6493E;
defparam prom_inst_0.INIT_RAM_05 = 256'h79F1B6FCBC2F207881398417A37CB04A52EC60828343E0C81E3B1A7DED9388A1;
defparam prom_inst_0.INIT_RAM_06 = 256'h80B0B0E14D90964808D8B03959297075ECF9CADE650F08ECA8BCA1DB6742DF56;
defparam prom_inst_0.INIT_RAM_07 = 256'h03377515D5393F2CBA791000BF209754BEDDDD27828A2084C1E02E828685A0A4;
defparam prom_inst_0.INIT_RAM_08 = 256'h37D94E689BDF3919594D45370038E8463E43C49252C22821880B07CBB8E24D1C;
defparam prom_inst_0.INIT_RAM_09 = 256'hE7F39B8E6B8E09512EB8EBDC073F15D6D1ED512B38D464850043DEF671666C19;
defparam prom_inst_0.INIT_RAM_0A = 256'hC75138161D3E8BB5DBED0538FBEBFC8258E288EF9B749CDCAB8A083405F6D090;
defparam prom_inst_0.INIT_RAM_0B = 256'hBBDC24EF8346875623B4689CE1D6A3D1273F45F05CC308BE47408475900281D2;
defparam prom_inst_0.INIT_RAM_0C = 256'hFDB044A7442071C9CAE090B1F54984B8C2CDF9D76438B95EA3085044108825EC;
defparam prom_inst_0.INIT_RAM_0D = 256'h65E49C092B080B27092B0801CAE0B3921541C939E72B82CAEFE786F344769736;
defparam prom_inst_0.INIT_RAM_0E = 256'h2E996A159F1554552C2C1D64E0759CF4609855979272B0B0A794A0C94855941D;
defparam prom_inst_0.INIT_RAM_0F = 256'hD3A095A59845389C8944279E694AA090838976C78C4EBC70A9C55495142A8E49;
defparam prom_inst_0.INIT_RAM_10 = 256'h7939C6CBED5EFDDE559FD279C63944E7FEEF12325D511527F9A43FE11279B19E;
defparam prom_inst_0.INIT_RAM_11 = 256'h1428E42E84414743EA3B90A3D49ED55CBD2792FB54A4A6608A4E49E739955552;
defparam prom_inst_0.INIT_RAM_12 = 256'hB495795954551D4F4F5797397C1CE39140ED1473800473781C738AF560883514;
defparam prom_inst_0.INIT_RAM_13 = 256'h4A98BD2D1925A49364D25A4996496F865C64F60900440930B5E2794A949C5546;
defparam prom_inst_0.INIT_RAM_14 = 256'h2ADC970EB43A095F574569A7519D49E51976702A12751A32C6F3B13BF592ED42;
defparam prom_inst_0.INIT_RAM_15 = 256'h954A2D2D420D0AD89DC504D29DCE5F45CA646AD32E2A277A07A126A72A145BC6;
defparam prom_inst_0.INIT_RAM_16 = 256'h75572B82B372D7F070F564671F24B3FB3E49C27DC78242426528B4AD08342750;
defparam prom_inst_0.INIT_RAM_17 = 256'h0BD28FE0BDEE3DCBBF20F21D5F275E1CC2623E352772FF13E195115656277619;
defparam prom_inst_0.INIT_RAM_18 = 256'hF6528598AD3196AB4552756827073B355D48E8AC253E37A3274905450C97E8F2;
defparam prom_inst_0.INIT_RAM_19 = 256'hC3BC58F6CAA1CBBF2D58659391996B289290945BB36B490795919382092536B4;
defparam prom_inst_0.INIT_RAM_1A = 256'h185956EC175E6BA053A9C2B46D6B55AD0D39D505848C85C23515464ED11990A3;
defparam prom_inst_0.INIT_RAM_1B = 256'hE8D2D66DD2652B489DC4569BD11A12565A4634606358C1EFD11A5699CC7CB11A;
defparam prom_inst_0.INIT_RAM_1C = 256'h0B2B46FA10514C9751C9123FF852B561DC61451C27848FFEF71C50741C0E14AD;
defparam prom_inst_0.INIT_RAM_1D = 256'hC7FAF85DA343FE5C7F24614B1D330BF2638161504B722B2FF0945547C9FC591F;
defparam prom_inst_0.INIT_RAM_1E = 256'h1CD96F4E51D12AF70AC9824E4271750792511D4D46510FB3FBFB2E2C3F3B7F28;
defparam prom_inst_0.INIT_RAM_1F = 256'h1D142F5953BFC6C45D765E718DD5126ED3BA564EBD18E1294E59D4B4F7A93AF6;
defparam prom_inst_0.INIT_RAM_20 = 256'h770BD9CB5449976462F58D9F42EB422BE447655D48D1954514C5153B1A415025;
defparam prom_inst_0.INIT_RAM_21 = 256'h2FB7AD28E158A8E22522B36E290A0962B59D089DD4AD539395D173D61A4B2523;
defparam prom_inst_0.INIT_RAM_22 = 256'h9582DC9D61A491452827888E57CA1717574A1D5D464AADAD55EFF3811A15D443;
defparam prom_inst_0.INIT_RAM_23 = 256'h41383435F1C636783AE000DEBED3834352DED46E409A9381D2F477C64A4A5551;
defparam prom_inst_0.INIT_RAM_24 = 256'h5996519D08E1886386CB61B238ECEF1C574E272591BDE8A28128341CEF1C1B42;
defparam prom_inst_0.INIT_RAM_25 = 256'h69C99D0B9665C8D06D6474619325D18236237DC65287599CAD251DD99B674490;
defparam prom_inst_0.INIT_RAM_26 = 256'hC104D47181B028DB499EAD1D259C9D4C9DE8ADAD66F612853A1C4142A48D9DB9;
defparam prom_inst_0.INIT_RAM_27 = 256'h7F0707291B63C265A5BCB076D52C1FBB01BE7278384966B81C1C06F239DE9152;
defparam prom_inst_0.INIT_RAM_28 = 256'h958460469442C1F1460BC4D6B762479EE798B072749257904692544C33462C26;
defparam prom_inst_0.INIT_RAM_29 = 256'h4693C095133F383165BE0C935A9CF04697643D04690607072E12490CD90B87E3;
defparam prom_inst_0.INIT_RAM_2A = 256'h551461946719571877F04800E5D894E7214C2E9391C112E924564901C1CA5630;
defparam prom_inst_0.INIT_RAM_2B = 256'h587B865C83C65F819AD0AD0211321B04493744C12B6FDC7187C6D4E654F7FF40;
defparam prom_inst_0.INIT_RAM_2C = 256'hDFEDD4D9FBA8D5471A1754567579DAD08D9DAD32ED622196FF8D193BF8EB8BAD;
defparam prom_inst_0.INIT_RAM_2D = 256'h37B9471F9075E5C34ED71D50894638E186CB39867D1D7E5CE6EC2ADC1DD275C1;
defparam prom_inst_0.INIT_RAM_2E = 256'h83B54A4879FA6E1355BF5C20E0EEFD3B84E477B92C1FBE0A154F752A1E7BF4E5;
defparam prom_inst_0.INIT_RAM_2F = 256'h4A6A39AD37464209037BB854559E7859619C3468DAD859AD74A4F41744CA2A18;
defparam prom_inst_0.INIT_RAM_30 = 256'h774E9DFE144A77C14A447415D054E393A2B7159919F89792709027820EC01E44;
defparam prom_inst_0.INIT_RAM_31 = 256'hBCBEB36383C627394E71512614E734E5BFFCA507786C9B145E49CEB8BDB36376;
defparam prom_inst_0.INIT_RAM_32 = 256'h0D144543979D4A2298A808D8BD8A0E9D06075F4640743DF8BD6567DB9457A234;
defparam prom_inst_0.INIT_RAM_33 = 256'hB19455E1FDF155D49D7BBE32FA8177B0FC29771B1C38294A189B70F121BF5EC2;
defparam prom_inst_0.INIT_RAM_34 = 256'hCA5505997DCFFDE022700019CCCD55D59A6716412DB90E403D67290419746271;
defparam prom_inst_0.INIT_RAM_35 = 256'h22C60A83FFF1703FF5D60E5AED578A05C8ECBE0359DCE49175707624F089207A;
defparam prom_inst_0.INIT_RAM_36 = 256'hB4E31729D7592140B790B82C661CAA7DE72A18B291B74293B7677CF2F22F292E;
defparam prom_inst_0.INIT_RAM_37 = 256'hBCAA1B511B074C997A4B1B1B7BB1DB89B221845FC0AF34099C0B1DC61B903292;
defparam prom_inst_0.INIT_RAM_38 = 256'h089D1039496EB02994D4E7925462DF85D11D275870BD039257B82F872746FDDC;
defparam prom_inst_0.INIT_RAM_39 = 256'hF85CB845343110A069F19EF728156B7117AAE1463B9478254AD9D0274DF274DD;
defparam prom_inst_0.INIT_RAM_3A = 256'h9B0F02D11D6475E1B138A18919B19BF186B4ADE568D26EC2B44631F98E49D1B7;
defparam prom_inst_0.INIT_RAM_3B = 256'h0A38ED113771C0F62873BFBB934219238C2F2C62AF405D4945BB2DB8CAC2A742;
defparam prom_inst_0.INIT_RAM_3C = 256'h565692808249429292D0D04953B65257E15C93E08DC45E50B04A4E3B24D78649;
defparam prom_inst_0.INIT_RAM_3D = 256'h51D51DF195C757A52B789C2095246755C63D4B4125C941B6C4671559518455A5;
defparam prom_inst_0.INIT_RAM_3E = 256'h0B9D42E059D9E9117BA3BE67627741013A5B5BD1DFF2A554D411F89C41E1181B;
defparam prom_inst_0.INIT_RAM_3F = 256'h0B76F46C271C2505DE7D56446A39147928994D4EE1BC60F0ABE527F82F28506C;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[29:0],dout[3:2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 2;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h0EFC3E7081F25FFFD4FB1F2800F51C1F83A571C9FFC8FD870FFEFFD02F3E23CC;
defparam prom_inst_1.INIT_RAM_01 = 256'hE1F484407A500D00789FD00C31338DF15C7105051D407B3619B9CEF109CBB8EF;
defparam prom_inst_1.INIT_RAM_02 = 256'h12F7835C5D05E66083440B9C20526154704F034D015F4CD4345453765EFFFDC3;
defparam prom_inst_1.INIT_RAM_03 = 256'h1501C41319AF7050D1F1E06C6744174B4F5384374D374E579F053174D104510D;
defparam prom_inst_1.INIT_RAM_04 = 256'hDCD2FEFEEF8EA95769B75FFAFB9EF88058F503BD44003212FE52AC456D55A233;
defparam prom_inst_1.INIT_RAM_05 = 256'hDF1E851EE939BD2EF00FCF4F4244EC03EB6ABAEE62D323A477B7BF3CFE04AC92;
defparam prom_inst_1.INIT_RAM_06 = 256'h6452CA8483B8E5844CBAA6222E110922D23BEBA784282C784AC7A114B2F840D1;
defparam prom_inst_1.INIT_RAM_07 = 256'hF413ABFBBA8A1B70C47F3D027F9EAC0C71FBB23BC3631402A6F91563AB02D95A;
defparam prom_inst_1.INIT_RAM_08 = 256'h2B5246902B128A0EDEE054341130BDE035271D771D8D65C5360C4B64CC7C2C5E;
defparam prom_inst_1.INIT_RAM_09 = 256'h253ACCC5FCCD61535FCC4CB2E0BB05CBAB88D0E9E9B4195A0391E2CBBA1FA060;
defparam prom_inst_1.INIT_RAM_0A = 256'h84E1EC52173C47E5CCF198F2BEFCFE7A6C9738FBC4E51BDCDCC14CA9B5137CFE;
defparam prom_inst_1.INIT_RAM_0B = 256'h57E218FBE5CDC5E3E09F605AB1331A333D8F8CB87C4B847385D1E45E4109D13D;
defparam prom_inst_1.INIT_RAM_0C = 256'h27CA4F836F6022A37A3DA1F381C8A2F076C2B48F1F00E4D4C9D80E4FFD076272;
defparam prom_inst_1.INIT_RAM_0D = 256'hFBBF35B7E9DBBFCFB7E9DB0B7A3DB3FB7DC0B727BDE8F6CB62BD8B61F223CCDF;
defparam prom_inst_1.INIT_RAM_0E = 256'h3074FC0D7701EC0627687DCFADE7372FA07CF3EEFCDE1D98DEFAB6078CF3EF38;
defparam prom_inst_1.INIT_RAM_0F = 256'h413D8DDFF4730CF663E7DEF9EF663ABDB8CF1F0A47038C83E6C073B608770FCF;
defparam prom_inst_1.INIT_RAM_10 = 256'hEFF3BAA0F4D0004177F01DEFBAFBAFCC0B989F93CDF6128DA7BFA011DDEFB97F;
defparam prom_inst_1.INIT_RAM_11 = 256'hA63FA63F2BF8AE62B80CA07CB23F4D4851DEF83D309F0FE07DF887FCFB5D49DD;
defparam prom_inst_1.INIT_RAM_12 = 256'h2FB834FD8AD0397EF0C05C85E6932F2B6BEABAEF206BDE3C82114E0500C4A2B6;
defparam prom_inst_1.INIT_RAM_13 = 256'hA7A0E321632800140232800137CB070F98B0040D9341104103FDEFC44D3C075F;
defparam prom_inst_1.INIT_RAM_14 = 256'hF242B2BC93BE87E8F8773F32EC09CC5DCB8342B3632C23C6BFF1061E06E1E84B;
defparam prom_inst_1.INIT_RAM_15 = 256'h13B4C3E3B4E384B8CB9E87B34B6DC8FE363F44B5FE1D32F1E3E6027DFA392032;
defparam prom_inst_1.INIT_RAM_16 = 256'hA2AB16036E2DB60CEBAD585A31707AF7ABF06C23AD43E3B27EDBAE4BDBAD32EC;
defparam prom_inst_1.INIT_RAM_17 = 256'hA5BB065A5B8BFB647FDAC3A30AF2D83128B2A72DB2DBFF4BDC94DDA3F5B2F70F;
defparam prom_inst_1.INIT_RAM_18 = 256'hED33AFF64B28FC12E7832E1A328E8EE6264E3A32B112EF6ED2CEB344605970E9;
defparam prom_inst_1.INIT_RAM_19 = 256'hFF00880087A0647FFB4D1FFF0C04FEBC48D8E5EEEE32FBE34FDC9FBC2D07792F;
defparam prom_inst_1.INIT_RAM_1A = 256'h0DC7FDBBCFE75FC30F3F592FEE12FB4BEBF05C8CCE52F879E1BF727E5724723F;
defparam prom_inst_1.INIT_RAM_1B = 256'h5B21C33B591D92E0CB82007024CB79FD3FDD2FC02906C80064C93F0748D8D9FA;
defparam prom_inst_1.INIT_RAM_1C = 256'hE892FE23BCC44679030771BFD65BED13AC3BCC48994C6FF56B08F02A0B2596FB;
defparam prom_inst_1.INIT_RAM_1D = 256'hDD81CEE0F2F05D7828783766039167F1E174375004919B1FD2EDAAA247FF8C39;
defparam prom_inst_1.INIT_RAM_1E = 256'h8005D6FA57D73B6CE740A3E70B780723F157F34C7EA308A3AA2293389AFFE87A;
defparam prom_inst_1.INIT_RAM_1F = 256'hAFE236E5CE003ADE7DE13F4C87DF621311897BC4DBE9F126BA6EE07B8C13E96E;
defparam prom_inst_1.INIT_RAM_20 = 256'hF0ADB40D7BF85EBFA36E6A34035883188D608C768CBF005D7A000EE0BF60F81F;
defparam prom_inst_1.INIT_RAM_21 = 256'h3D5BCB107C36FE7BE2287B161F0C0CF72DCBEACB4DCB817E2783701E0FC71C92;
defparam prom_inst_1.INIT_RAM_22 = 256'h002EBC71E0FC689D3C1E463AFE3A8EBE1D72F3447E7ACBCBFE400F88F98C0F0A;
defparam prom_inst_1.INIT_RAM_23 = 256'hA6E38F4E892508D8E180007FC76EBAF6ECBF20F3AC4FECACBB6FADB285F03B4F;
defparam prom_inst_1.INIT_RAM_24 = 256'h149D7E10E3CF2F4C3004DE01E3034A38473CD2E37F2AB72D30C38C0B82B88F34;
defparam prom_inst_1.INIT_RAM_25 = 256'h27C7CBF37BFFD4B2FDC2AFCEBB1C7E892C32E7FD334D7076CBED8FB07FF2CCCC;
defparam prom_inst_1.INIT_RAM_26 = 256'hB4C00DC1DAEBE87AC7F6EBDBED4FB024DF52B4CBFF6D3D00E175C07EBDCBCB6B;
defparam prom_inst_1.INIT_RAM_27 = 256'h4D1799315183D04DF5007178F71C5DF1120047747C7081345E6467B0CCBE7B8B;
defparam prom_inst_1.INIT_RAM_28 = 256'hDCC791B1E111C5C4441F0C84080384D3F5C0717055E77501B1E7751034791C74;
defparam prom_inst_1.INIT_RAM_29 = 256'hB1E4F1DD447D3C370C1C0DE2101FC1B1E4953E1B1E6717990D538E0D1EC34FC3;
defparam prom_inst_1.INIT_RAM_2A = 256'hE2BAD2F84DC952FB8C000D72011023380A0CCC11E4F104C105700545E64DC441;
defparam prom_inst_1.INIT_RAM_2B = 256'h87E4F260E83267A97CB4CB01002103059170598A4008882EAEB21301772E0068;
defparam prom_inst_1.INIT_RAM_2C = 256'h008A982344FF85AED973740B2FCCB4B64BCB4B201AB11F73004BC2FA7024F756;
defparam prom_inst_1.INIT_RAM_2D = 256'h024E51A800137E60A724EB8E3074CB0CB004E37A88C3017B2B141DC82A34D0A3;
defparam prom_inst_1.INIT_RAM_2E = 256'h88688707D8F67C0A3601FC363ABB02FA627E3A4E1F045C8F78006A1DF52C0BE6;
defparam prom_inst_1.INIT_RAM_2F = 256'hC1CC8E4B8E2BFEF3BCEC6E8AD2F0E02F4A37EFA4B4BDC74BFC1FCCA1428C9D8C;
defparam prom_inst_1.INIT_RAM_30 = 256'h2D664B02B40FCC806D8FAC82FF16B37E992D9CEFE276EEFFCB7ACD4F6BD83D14;
defparam prom_inst_1.INIT_RAM_31 = 256'hEA6BEE1859B20DEABC172715C3CEE7EAC000F829E6F27E8E3F437E62DB6E12E5;
defparam prom_inst_1.INIT_RAM_32 = 256'h6AB48CDC994B387E983E64B4DBCB6B4BE30EDC2CFBBE9A20DB17BC94E234CB2F;
defparam prom_inst_1.INIT_RAM_33 = 256'h2EA0D8973E79BEAD3484C1A313013996E63D943F892DAF03F27C94993F00AB0B;
defparam prom_inst_1.INIT_RAM_34 = 256'h44CD7B38CAD5D8D63F3AAA901DF881FEB7AFCAF839C5AF80AD54EA81B3EF4C1F;
defparam prom_inst_1.INIT_RAM_35 = 256'h2DC44789554188AA95E7C06C35F784CB8F3CF3099C0487127DE1C5DDC3CF1C67;
defparam prom_inst_1.INIT_RAM_36 = 256'hADCB79E2E76E1C30F60D0F62BA8FAD9D92AEBC7EB77D2E3D3AF2D04242E42515;
defparam prom_inst_1.INIT_RAM_37 = 256'h8AAEBF0137AADAB379CDF2D0A4CD3C4CF13DA4CFE8741ADAF2DAEBB2D3C6EC83;
defparam prom_inst_1.INIT_RAM_38 = 256'h3F3684F663ACA41871B7AAFDCBCC3970853F12E738DB8178E64F6AF3FF13A6BF;
defparam prom_inst_1.INIT_RAM_39 = 256'h89BA3A4CBA393CB6F5383D6D9F0FD2C939E77C3CFAF3C763D4BCB692DBB12DB6;
defparam prom_inst_1.INIT_RAM_3A = 256'h0DA4A148D3DF6D3F97DB0DA73B07702D8EE20D17F6613BB8BE0038EF6BF363E8;
defparam prom_inst_1.INIT_RAM_3B = 256'hBFDBCE93FD9A64401033C244E33ABB830F83BBEF36C82B44D94CC3C4472AF3B4;
defparam prom_inst_1.INIT_RAM_3C = 256'hAF7A3C30F18EF97FAD3EB42EED2BE3BA00B5D9B7DB84EBEBF2C5FED3DC7F0DDE;
defparam prom_inst_1.INIT_RAM_3D = 256'hDF35DB0772BCDAD0C270376832036EE7BAEB72D0BB2DC0DEE2CCB78ED726DE37;
defparam prom_inst_1.INIT_RAM_3E = 256'h2D4B4753F4BE3D93BEFBEFB2FB2C0CB8A7B75C1F38ABE02DDC010E3280AAD84D;
defparam prom_inst_1.INIT_RAM_3F = 256'h3F9FCEB23FFA3F87EBFFFD14CC8E84EFE04F1B7A73D0B243F417126076E3F2B7;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[29:0],dout[5:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 2;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'h6CD6962E8BDEBFFFD07E3E8F84C43CBDE9EB5268FFF4FF4C4CD6FFDC159643DB;
defparam prom_inst_2.INIT_RAM_01 = 256'h01090955400500554140110101401001008105152011404064001C5B8DE775C3;
defparam prom_inst_2.INIT_RAM_02 = 256'h540414511051040410111000410104410A1028104410410402011440403FFC04;
defparam prom_inst_2.INIT_RAM_03 = 256'h5450044400400111150505015014505000540580604010041010410114440051;
defparam prom_inst_2.INIT_RAM_04 = 256'h8CCBAEA403A0000057577D5AB7F57CF8AFBA3EFFA21F495F010F001F411F4140;
defparam prom_inst_2.INIT_RAM_05 = 256'hC3B4E3B4C8B2B4AAD244AD2FCAE2C480075C72CFB0B97F04789AEF3DA25521C8;
defparam prom_inst_2.INIT_RAM_06 = 256'h024FDA0661C7C82007324E028D108828020CBFCF42309DBC49ED338E20D3E321;
defparam prom_inst_2.INIT_RAM_07 = 256'hAC2E39094CBCA03584338000C0E4C46402B33C31CB2B5A3A002002EFEF38C0D0;
defparam prom_inst_2.INIT_RAM_08 = 256'h5154E40500313D650533F01438AB353C2CF2F30280F130A2F36E6D7226B5B235;
defparam prom_inst_2.INIT_RAM_09 = 256'hF0230DDC3DD81E3A82DD0F9418B128E30CAB264C7EC1F2D801120EC33CF60580;
defparam prom_inst_2.INIT_RAM_0A = 256'hB23BED1BC830E9D8ED3D1303DDFD0393CDC33D77F251138ACDD03DCF6233AC92;
defparam prom_inst_2.INIT_RAM_0B = 256'hC8BEA977C2EDD203CBEB07133482C1923451C904D3217082D23DF7203ABCEC84;
defparam prom_inst_2.INIT_RAM_0C = 256'h8DE6B1006DF08F2C9037CADEAA402F029F303EB33756C25E0A7C4EB107E5FCF4;
defparam prom_inst_2.INIT_RAM_0D = 256'h54610858427CAD4058427CA09037CAC4D3424D0D6240DF6B12626BA372C33637;
defparam prom_inst_2.INIT_RAM_0E = 256'h01F43FE44E164448C9F9D359234D6D5960D34D51842427D43582310DA34D50D3;
defparam prom_inst_2.INIT_RAM_0F = 256'h8B37E62492F98CD2B62F145E798C3037C8CD93ECD42B50CBC1F99000173C2B4D;
defparam prom_inst_2.INIT_RAM_10 = 256'h41599680FE6BB9F94FD00041965961640889BFA3640104DBB9E4654BE145444F;
defparam prom_inst_2.INIT_RAM_11 = 256'hBA3D28339226728E74AD58B5680FE698F004103F943D2248B252110659508600;
defparam prom_inst_2.INIT_RAM_12 = 256'h0C02643E1612E915959250652309659C4169872586123E7E61BD2D695AEB61C0;
defparam prom_inst_2.INIT_RAM_13 = 256'hB316C0BEF0BEFAEEBA0BEFAEAC2EBAD2EAEAFBEABABBBED009F145DF24085952;
defparam prom_inst_2.INIT_RAM_14 = 256'h4C112453067D5BF004048000C5F22C7F5C480B70080DBB1555475650095142B7;
defparam prom_inst_2.INIT_RAM_15 = 256'h8F124242124220360320E4CB0346C03101FC4030D55D80C035C2A57D48034ED6;
defparam prom_inst_2.INIT_RAM_16 = 256'hE0AA202B07A7200105C843938B0F94094316154030B7F3120C490803490980C4;
defparam prom_inst_2.INIT_RAM_17 = 256'h293E2422D3AB469C80E44B082100EBB971A92CCC80E3150DC5E111F40480C0AF;
defparam prom_inst_2.INIT_RAM_18 = 256'hF9036676831FF000F4500C15BEEFACEC556D3D3237C5339300ECC0C518A3228E;
defparam prom_inst_2.INIT_RAM_19 = 256'hEAEC0D9DA0599C80C420CCC4A5F43FAECACAD51847A0C03643F5E4935C9F020D;
defparam prom_inst_2.INIT_RAM_1A = 256'h20330021E20E68C9648B880D2800C403424A7EAF0133D2FC6BC0969202573330;
defparam prom_inst_2.INIT_RAM_1B = 256'h41115B0405CC80F6034981FECD5804010F10CDE0A58FD9BB8D590F3FDE3A044D;
defparam prom_inst_2.INIT_RAM_1C = 256'h4C80D368060AA3B41E4D40C00B80100E9E8020A6E038300227ABB227A8B2E004;
defparam prom_inst_2.INIT_RAM_1D = 256'h51D24F120CF6C8F4BD3D0C012C6639E8C8BA0C20B3236EA015C0AAAA9F0320E3;
defparam prom_inst_2.INIT_RAM_1E = 256'h7B8500D6545453CC3740F7B3F78ECC0B71D47E9E9E28DDFDD444098BCD013D33;
defparam prom_inst_2.INIT_RAM_1F = 256'h5048ACC525AA963D43E90FA594400088A53D4614B3493F68169518515954580C;
defparam prom_inst_2.INIT_RAM_20 = 256'hC0AF340D4512526122CCB82A205627E6A012594CCC37AA514600705A0F17153E;
defparam prom_inst_2.INIT_RAM_21 = 256'h70834332F48531E368A51C20CEDDEF220F834C83944320F598948C316DC73EAC;
defparam prom_inst_2.INIT_RAM_22 = 256'hA9146CF316DC6531B75F2B530292627253927E9A9E92834300FBA4994C517F24;
defparam prom_inst_2.INIT_RAM_23 = 256'h6179D9C9BB2CE5AEE3A0002FD3179D9C976FCE3B6003C69662CD5A9A0BD28447;
defparam prom_inst_2.INIT_RAM_24 = 256'h523CF48A4D34FDA69A8E35A349696AE846527B7B67ABBDE7B279C809EAE88E5E;
defparam prom_inst_2.INIT_RAM_25 = 256'h0FCFC34C77208332354F7165973D858ACDB0D421037143F18301D883F100F805;
defparam prom_inst_2.INIT_RAM_26 = 256'h127403C9C8DB7D450037D44201D80576D803338322CDC5824AFFC2F7C03383D0;
defparam prom_inst_2.INIT_RAM_27 = 256'h50BEBB8546AABBAB2AEEABCFAAAAF2AFBEEEDAEAEAAAB942FAEE5001843CFE0B;
defparam prom_inst_2.INIT_RAM_28 = 256'h2AAAAAAB810AAF3EBB902A01010AABAE8AAEABEBAB8EAEEAAB8EABBE45AAAAA0;
defparam prom_inst_2.INIT_RAM_29 = 256'hAB8FABAAEDAAAA441AEBEBA804FAAAAB8ABA88AAB850BEBB90542A916AAEAABA;
defparam prom_inst_2.INIT_RAM_2A = 256'hF187098A9B6A5A5909401ECABAE6EAA9BFEEBBEAAAAAE7BEBBAB902FAEE0ABFA;
defparam prom_inst_2.INIT_RAM_2B = 256'h66265693469690E5843283100000041435014318D8FBBB24BA9A4169455A002B;
defparam prom_inst_2.INIT_RAM_2C = 256'h9BB89396A64D2B3A698908000C003031B383031542515468AAB3594942F65A40;
defparam prom_inst_2.INIT_RAM_2D = 256'hEE2050DA901050FACB985626969A69A69A8E58D628622949A19E2D180901ADAB;
defparam prom_inst_2.INIT_RAM_2E = 256'h110800F51E1900BEC8ED4272723BA84A6F532220016010DD4211080145A2A128;
defparam prom_inst_2.INIT_RAM_2F = 256'h03CC4C8372261A6A59A663070189A0586D69992330303303213DF9496F144444;
defparam prom_inst_2.INIT_RAM_30 = 256'h0D2B03A9810FBD012D410A650698A876FA0D50584ABB51850581422B2F5EC50B;
defparam prom_inst_2.INIT_RAM_31 = 256'h4243479408131A58529F8C35592CC924EAA831972239CE610F269642B3479CE4;
defparam prom_inst_2.INIT_RAM_32 = 256'hD9C14055A143DB26F2B16736B32FA343BBF918ECBF21ECECB39462A64504C9CF;
defparam prom_inst_2.INIT_RAM_33 = 256'hA58B96980B2C50906922287F943034C6873E368D808CBC2B59CE22E105AA3B8F;
defparam prom_inst_2.INIT_RAM_34 = 256'h80C5102D890F58D4EA35555578F3198D8C6346349A651DAACA504478E8B1A5A5;
defparam prom_inst_2.INIT_RAM_35 = 256'h086241C000280C001C4088041861C24086144101C61C72081060400C61860701;
defparam prom_inst_2.INIT_RAM_36 = 256'h0D0D42434180048EC147ADE1012111E27ABF8C14CF7217F4E730D45050850607;
defparam prom_inst_2.INIT_RAM_37 = 256'h063F8D02C424160F73C55A5A66646640E2358B0C2CB0A64D8D4D569A4BE6C4BB;
defparam prom_inst_2.INIT_RAM_38 = 256'hAD0A76DFEC2CCA287ECDF18501272BDEB2C8B0E4063333FB0221E983503CC811;
defparam prom_inst_2.INIT_RAM_39 = 256'h778B22B003A2C6F23016874FFD6000DAC3AA3592498B15FC003C3D30EC030EC8;
defparam prom_inst_2.INIT_RAM_3A = 256'h4E98BB9C524148D5924D24B354E47EE4B82B0A940300339AB3202E98161088D8;
defparam prom_inst_2.INIT_RAM_3B = 256'hAF5966AC523CB0C03AA072A6505A54C0A9A9B1260CE5100602224220CB9BF413;
defparam prom_inst_2.INIT_RAM_3C = 256'h3900F4AFF1A50776872722F505A6294401E2F662EC2B060AD30BD65950C03424;
defparam prom_inst_2.INIT_RAM_3D = 256'h17E842E8B69F8EF17A4369E36535A21896461C8BD414006003A0643532279010;
defparam prom_inst_2.INIT_RAM_3E = 256'hAEC32B9E0C370CAC1DF5DF20EA0C2ECBCD409707EACBF600400109E3468C6846;
defparam prom_inst_2.INIT_RAM_3F = 256'hAD1340BE81CE80A04614010B0C4E2B18408BECDF8BE6B98ACE9402A2BA460ABB;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[29:0],dout[7:6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 2;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'hCF54147FC258FFFFCF471DFFFCBF4C25414F2F53FFC7FF07C754FFCF45143FCB;
defparam prom_inst_3.INIT_RAM_01 = 256'hD759595D77575D75D75DD75D75D75D75D595D7756555D57765575B5000CC3CF3;
defparam prom_inst_3.INIT_RAM_02 = 256'h755D55D757555D55D5755D75575755755855615755D5D55D745757757562235D;
defparam prom_inst_3.INIT_RAM_03 = 256'h55755D5D775555D5D75755D5D5D575D5D5D5751745D75D755575575D55757575;
defparam prom_inst_3.INIT_RAM_04 = 256'h33300027FC300000DEDDE7FAAD67DBAFBAAAEAAAFF5041505150555055505757;
defparam prom_inst_3.INIT_RAM_05 = 256'hC71400177C1C243090C3C90700007432F3573CF1C33170CF140C7F3C0EFFEF37;
defparam prom_inst_3.INIT_RAM_06 = 256'hF0C0F1C402CCFBCF34F07C7034000033701C037100DC0F341C450C00F3D070F1;
defparam prom_inst_3.INIT_RAM_07 = 256'h70C3FF1F14241D7CCF030000C0350CCC130CDF4D33033801F33CB3838303FC3C;
defparam prom_inst_3.INIT_RAM_08 = 256'h883258A3232CE572F2C100A58CF032C0F6C32C3133C33070CD484A1444960232;
defparam prom_inst_3.INIT_RAM_09 = 256'h90D00FC00FC03C3083FC4330201C8C0FCC53FF2E40F0D8C6019265D87288B721;
defparam prom_inst_3.INIT_RAM_0A = 256'hC3F24C030FE4CCFC0F0C0F30CF4F00D4FC03C73D00C0CC8C0FC40C7710C06470;
defparam prom_inst_3.INIT_RAM_0B = 256'hCD1C3B3D32C033F372593E0ECCF0803E1C0478C07000201373F3DC3F30CB30F8;
defparam prom_inst_3.INIT_RAM_0C = 256'h07400CB3014003CBCB3513FBCFC0093094003C3F0F0003FC0250000CB53D4F3C;
defparam prom_inst_3.INIT_RAM_0D = 256'hCB3CBC0F2E500F2C0F2E5007CB3512D071D003033F2CD40B1F3FC3F1C0701C1D;
defparam prom_inst_3.INIT_RAM_0E = 256'h8130F33C7203CC0C794C71DD41C7715D4031C72CF2F2E5020CF0F40351C72C71;
defparam prom_inst_3.INIT_RAM_0F = 256'h80353F1C709C0C7007091C7DF7CB30C500C7F087CC02064040F3FC3CCC3C0EC7;
defparam prom_inst_3.INIT_RAM_10 = 256'hC75314C3C3F113707F7031C714533D4C01102421F0D4001CF7DC300271C73C7C;
defparam prom_inst_3.INIT_RAM_11 = 256'h20B54FB5C0F32FC0200803D57C3C3FFE331C70F0FC0D41C3D1D4071C531FF3F1;
defparam prom_inst_3.INIT_RAM_12 = 256'h3C3220F3F3FFBFD5D5FC1C01C03D450BC14CF2F500C0C3F330F0080FC2FF3CBC;
defparam prom_inst_3.INIT_RAM_13 = 256'h433CC3855485545555485545552155525454554550551558FFC1C7C43CF80F3F;
defparam prom_inst_3.INIT_RAM_14 = 256'h4080101021010C10CF0703D3F631C04F60F00200013C2015555454143C404043;
defparam prom_inst_3.INIT_RAM_15 = 256'h17D86767D86704F04F0FC030CF7320D3CB2C74F10B8013D30814033540B33454;
defparam prom_inst_3.INIT_RAM_16 = 256'h7C010F03B4347C30C15F30BF010BE34E30D846030D0B0BD85F619F4F619C13F6;
defparam prom_inst_3.INIT_RAM_17 = 256'h05F307F05FA9675CC0706030F3D3CF0000A8333C13E06000C63F1F9CFC13D000;
defparam prom_inst_3.INIT_RAM_18 = 256'h1C3040704FC0B0D3DCCD3F733FC3073FFFC337B07F200DC0D3C007C80C3D307F;
defparam prom_inst_3.INIT_RAM_19 = 256'h9556FC04C11C5CC04BC01CF63630F01CD3D0F3FBF433C3320F36361881133E3D;
defparam prom_inst_3.INIT_RAM_1A = 256'hC1C71FED02F678418607413D8BF3CF8F67635FC30C0098455347D8D877CCB833;
defparam prom_inst_3.INIT_RAM_1B = 256'h03C060CB732C13D04F4001344C50701C3C2E3D40000C08118C503C03CC100061;
defparam prom_inst_3.INIT_RAM_1C = 256'h5013D814BC33C7C00B0140500DF02F0BCF0BC33CF02C140373CEC033CC137C0B;
defparam prom_inst_3.INIT_RAM_1D = 256'h1DF38D3C23F059743F0CCFC10C31BE1340D3CFF423D735F0183500175C01C3B1;
defparam prom_inst_3.INIT_RAM_1E = 256'h1131E3D4CF4F0D3C0340030303C0CB3370CF47C4D0F0CF70F333010CEF33FF00;
defparam prom_inst_3.INIT_RAM_1F = 256'h035013F0F500140C70CC3CF50B0D401132E4B1CB4F53D654D4C4201D5C07523C;
defparam prom_inst_3.INIT_RAM_20 = 256'hCB84F0C0B0D42F1D4D3FCC78033003F055FC1CB3F4F43F3CF3C00F50CD00C00D;
defparam prom_inst_3.INIT_RAM_21 = 256'h04DECF00650F30605000C5340C0D0F1D3F8F434F834FF0350F0BC32C8DC30E13;
defparam prom_inst_3.INIT_RAM_22 = 256'h3F067C32C8DC333F006D00981FD83F1F2CD847C4D0D88F8F1F1105084000DC07;
defparam prom_inst_3.INIT_RAM_23 = 256'h03511D9F300001EC80500070F07511D9F67CFC313C0375357D3D5E14C0D8CFF4;
defparam prom_inst_3.INIT_RAM_24 = 256'h0CCF34005186014514200508514143BC021463437403018400611C4143BC8218;
defparam prom_inst_3.INIT_RAM_25 = 256'h03C3CF61B01CB4FC3C793D45330CB5113C13C30C302CB030CF0C087033F3EC04;
defparam prom_inst_3.INIT_RAM_26 = 256'hD45000C0C0C040B0C07C03570C08321C0F3037CF1E3CB4004071C0C40F4F8F4B;
defparam prom_inst_3.INIT_RAM_27 = 256'h55155515575151557554515D5514575515555D54545555D4555455D8B8FC3B01;
defparam prom_inst_3.INIT_RAM_28 = 256'h754551555D51457555154055755145555D545151555D5551555D555455D51457;
defparam prom_inst_3.INIT_RAM_29 = 256'h555D515555D514555D55455155D551555D55111555D5155515D5451575454551;
defparam prom_inst_3.INIT_RAM_2A = 256'h1CF2C075DC5313515C30035155545555000635515551575515555D455545D551;
defparam prom_inst_3.INIT_RAM_2B = 256'hF0F454F80014F3CCFCF04F000000039334C93348CBD111F52C143D4C7D5C00C2;
defparam prom_inst_3.INIT_RAM_2C = 256'h311CF0C7B4414FEF507C3C0F3C78F8F0CF8FCF044710CF01008F50503094513B;
defparam prom_inst_3.INIT_RAM_2D = 256'h4744300EC0030F30B90F57F518D4514514205014CF57C0714D1CF48C3C15EFF0;
defparam prom_inst_3.INIT_RAM_2E = 256'h111F01C3C47CCC24FF447C70707D0053090C3C440500CC0CBF111C04F034014F;
defparam prom_inst_3.INIT_RAM_2F = 256'hC0C0038F0F01D45315C47032FC7DF307C0795D4CF8F1C7CF2C0D1E3DC9000000;
defparam prom_inst_3.INIT_RAM_30 = 256'h3F098F003FDD1CC0002D5F3C353FB1B5313F1C07514D2CF3C0F02F0303C07C30;
defparam prom_inst_3.INIT_RAM_31 = 256'hF074B401C0D4DE53D8D7CF0D618FBD8F40033FC0F030B73CF00794F04FB423FF;
defparam prom_inst_3.INIT_RAM_32 = 256'hCCBF2F553FCFD435303004F04F030F8F0300CFC1F020E7474FCB1CF47CFD013C;
defparam prom_inst_3.INIT_RAM_33 = 256'h053EF3C711473FC57B044031000003E07077C30F1C3C0C0350B4E0BC0500E139;
defparam prom_inst_3.INIT_RAM_34 = 256'h4004545111140119549AAAAAABAEFCF43C0F80F00F470C507BCF2CF00B0D4635;
defparam prom_inst_3.INIT_RAM_35 = 256'h0010804000000C000C308201003000C042041080C20820020C2000C000C30330;
defparam prom_inst_3.INIT_RAM_36 = 256'h3CC07F2EF3C40000DC4505401044BF77130D0C32C32F040523E3C82020020300;
defparam prom_inst_3.INIT_RAM_37 = 256'hB0CE0FFC3302C0C730C153503445744CEEC530FF07D520507050571453C07511;
defparam prom_inst_3.INIT_RAM_38 = 256'h0CBE302DCBCF70787CFD0CF1FD457D943C3813CB30CF0032FF454CFE3FA64440;
defparam prom_inst_3.INIT_RAM_39 = 256'h2CFC300F3CBC383030E0FE7DF581E3C03DAE161860F3CD4C78F4FCD3CF3D3CFC;
defparam prom_inst_3.INIT_RAM_3A = 256'h83CC23C3572D5FC517514507CF4074752C3C0F0700003D143C30F2CF03CBC3C3;
defparam prom_inst_3.INIT_RAM_3B = 256'h0D514C030FC380000FF31F444014CF0CFD401D40D3F3CBC3534457473D00D3D4;
defparam prom_inst_3.INIT_RAM_3C = 256'hDCBC7503D052C07535757092F501D4B2C0B7333CCF00F3F0F1C0D4531C7302F0;
defparam prom_inst_3.INIT_RAM_3D = 256'hF47F57307FD1FC0F633079807C0141CF1457D9C24B01C01CF02C0FF2F7003F0B;
defparam prom_inst_3.INIT_RAM_3E = 256'h0F8F03C0BCF0F003CFCCF4E3F13C024244B3F1F47F00DFF50C01C37004C05001;
defparam prom_inst_3.INIT_RAM_3F = 256'h2FF03F3C1CFC1C07F3CF1C30C003F0CF2DCBCFD0C0F03CC0C00703F03F2CB03C;

endmodule //Gowin_pROM_0
