//Copyright (C)2014-2025 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.11.03 Education
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9
//Device Version: C
//Created Time: Sun Sep 14 09:39:45 2025

module Gowin_pROM_1 (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [12:0] ad;

wire [29:0] prom_inst_0_dout_w;
wire [29:0] prom_inst_1_dout_w;
wire [29:0] prom_inst_2_dout_w;
wire [29:0] prom_inst_3_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[29:0],dout[1:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 2;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'hA1F7273E7505F53A3AC46083B6861B3E347B49DF4D0119737E97D27860AF7D15;
defparam prom_inst_0.INIT_RAM_01 = 256'h691BD35E150A9DBD374A6F29BF782C25B56B4218376C0E0DE45696656045E5A8;
defparam prom_inst_0.INIT_RAM_02 = 256'h42EEC554B55864A71C56771C97461D08D5946460BD3BEA4F5BEE823B2C5BB16D;
defparam prom_inst_0.INIT_RAM_03 = 256'h5674F862E3A0B19DEBFC6311F1B1460AC619189C72DA5271D3B06293959D3919;
defparam prom_inst_0.INIT_RAM_04 = 256'hACBC2ED3E2E2CBE1EE85C42CCB08DF8AB2FD3A0158AB2F069A0A9099EDE17DD2;
defparam prom_inst_0.INIT_RAM_05 = 256'h1C47E6D3A3A475797D4D938E9F5E7F38FDC23FFF18E42E8FFED0A10FD84D5280;
defparam prom_inst_0.INIT_RAM_06 = 256'hD1B6178612414531E1B8D2B028174527E3D0B4686F92728B78619575717C7FF2;
defparam prom_inst_0.INIT_RAM_07 = 256'h68B9AC6095C816A09D2C615A15956D14F2BC68524E56660F280727E49CFE60B0;
defparam prom_inst_0.INIT_RAM_08 = 256'h1D734F44A1F4461AE134F44A04E3D1187634ACE09C235C0144DD128734461D39;
defparam prom_inst_0.INIT_RAM_09 = 256'hD2EF15165D44470195C15CC31C0941CF581F54BF7461726355D14A08A1525548;
defparam prom_inst_0.INIT_RAM_0A = 256'hACC54162C5095CC6B3B600A54B2270BF544AF59D29B160B681CA29B056289859;
defparam prom_inst_0.INIT_RAM_0B = 256'hB411DFBCA637EE8BB35E2B82BB974471DC7417CFC9FE8E3D8BAC24ECB9C2FF7D;
defparam prom_inst_0.INIT_RAM_0C = 256'hC6434197F519EE9269C57DD8E70A9CBB376EC9BF0F04532CE2D64768040B3774;
defparam prom_inst_0.INIT_RAM_0D = 256'h22280812B8281C67731C08E60A242746C78ABE0DF11A761BEB949CDC441A01CE;
defparam prom_inst_0.INIT_RAM_0E = 256'hCB927551B8FB352899D0FFB44568B86CD42E099968875C83A72740B3F5E29E3B;
defparam prom_inst_0.INIT_RAM_0F = 256'h32FEFBB86CDCA64F0B341B82D12CA17446555E820B761D0A69CB7CFD78EC0702;
defparam prom_inst_0.INIT_RAM_10 = 256'h742D4637C469146DC2653572CDF0AAE1934754CF17587412340E35385949CE7D;
defparam prom_inst_0.INIT_RAM_11 = 256'h3B3F2411564630A778DE01C05D09C09FE4A179D61AFBCE464DF4ECE1B5E1B60D;
defparam prom_inst_0.INIT_RAM_12 = 256'h0D398DFFE10F37CABCA39A393343C07554342D38745501A2208A0BB541EF853A;
defparam prom_inst_0.INIT_RAM_13 = 256'hA55091B425D0606F8206706878702743D0BC187BF9FA7EEC8BC7F4D46F11DC1D;
defparam prom_inst_0.INIT_RAM_14 = 256'h38A64275195C2715741BD116740BA70B1B97ED61E958457B86FB1D87C561D21F;
defparam prom_inst_0.INIT_RAM_15 = 256'h9D85116EF54A9D53465611495746CDEFF19D59DC467548BF019FDD864D950677;
defparam prom_inst_0.INIT_RAM_16 = 256'h02F4B46C4989D09C54B794A18A20B286B4EB19FE5C6722C0534A42C82BC58BD1;
defparam prom_inst_0.INIT_RAM_17 = 256'h6BBBBB19C6F5C7C751A5C6FC6D7D586E4FF5E56FD451354613D219F7544B45D1;
defparam prom_inst_0.INIT_RAM_18 = 256'h452872FBC4DFF7E5C645765F217C602F85116287BDA1C549D45143965C112894;
defparam prom_inst_0.INIT_RAM_19 = 256'h72193BE1B1B33043C6721C329DE21DC29DCA7FB35A7E09B0509E3638D8DD41DC;
defparam prom_inst_0.INIT_RAM_1A = 256'hD2D1074116C01D4F437494E3D0130719435CE9C7C94B21D7A09F1816D65575C7;
defparam prom_inst_0.INIT_RAM_1B = 256'h524CF627224DC9D5DC1464C62CE9FFFD5F9CDDB52CFB4E352F5BD7DC9275BD6E;
defparam prom_inst_0.INIT_RAM_1C = 256'h6FF25B79E1D1381F95C22BDEF34F46551DDDD8282D5A8BC552D38E27738A6EDD;
defparam prom_inst_0.INIT_RAM_1D = 256'h5457F6FDE106D826756C9279CAD3925618ECD0CA147A0437B58527C07FE625BF;
defparam prom_inst_0.INIT_RAM_1E = 256'hB1FB6DB964870BA0D075ECD0FA3738206053D54B4611903A4F2B549915C47594;
defparam prom_inst_0.INIT_RAM_1F = 256'h5CB40463EDFB77618D5BB555BB6FBB67EE55432EFD454EEF329515544B6F2FA1;
defparam prom_inst_0.INIT_RAM_20 = 256'h25C3560DD7D39D51D75E474C3F7FD556D75FEFFF0BB76EEFEEDD8AC9D4410041;
defparam prom_inst_0.INIT_RAM_21 = 256'h075501ED559D3A1C57475F7558A7BB055C87378414257DD587C2ECBDCBBC7CFD;
defparam prom_inst_0.INIT_RAM_22 = 256'h5BF6FF86D24FE3FD9D0B911C1B600C1AFF7445770DD735CD7359544665673963;
defparam prom_inst_0.INIT_RAM_23 = 256'h168D9670D95C6590655375F0EC545E55501C01FB5D557EDFEF1574049C043C8C;
defparam prom_inst_0.INIT_RAM_24 = 256'h24333FD10A5663EFC0A002B52CBEEDB430BEF8E2CEE2FE1908A18E5D1534D15D;
defparam prom_inst_0.INIT_RAM_25 = 256'hDDDD41DDDDDD1C5C8F42E02B5040014EFF73705D8C2C39BFF753BA57E0FED3B3;
defparam prom_inst_0.INIT_RAM_26 = 256'h8EB2FF2F2DE475D3874C4C6DFA3EC5ABAA3156CC4088AE3F8CFBB61A4A4191DD;
defparam prom_inst_0.INIT_RAM_27 = 256'h1054E387D5D12F5A2B8E8FCA7575E47547711D5751571394B57D6E4ADF54F502;
defparam prom_inst_0.INIT_RAM_28 = 256'hFE23CE2058E4D9A7E7936062379DF3DBA65F1C90B5571F595797124254B7F857;
defparam prom_inst_0.INIT_RAM_29 = 256'h3815C52EEED5DF134F40BF44642416C4F555D953A5019559FEF1505567D1755F;
defparam prom_inst_0.INIT_RAM_2A = 256'hF44A4718D05C34755D5F0D7CF74150D4F216EF4C5E3317CCC5D7FFFFF27EF416;
defparam prom_inst_0.INIT_RAM_2B = 256'h3675BC51D7DD5F846B7A6715085557D18611461169D155D57554D115450DD73F;
defparam prom_inst_0.INIT_RAM_2C = 256'h4D57F54E44D5F95A6CC059951AE285E949CE655D979193B14064D9D18A26571B;
defparam prom_inst_0.INIT_RAM_2D = 256'hCC54F290E80F3DD88464B377F478474DC1325209D0C134635D5773FBD5FF95C1;
defparam prom_inst_0.INIT_RAM_2E = 256'h338A36BE08CD2B5CA045A413821EE439070750F4005C0D12887035D0B710B1D2;
defparam prom_inst_0.INIT_RAM_2F = 256'hD153FE1E57786AD447742DD56BF58FF22DD15FF83674E27520376777F92DA1D3;
defparam prom_inst_0.INIT_RAM_30 = 256'hFFFFFFFFF46563441A30705CA074FED3474F45D30D4B81F9A58B0C624C446E0D;
defparam prom_inst_0.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3A = 256'h002000000200000002000200000000000000220028082A200820000000000000;
defparam prom_inst_0.INIT_RAM_3B = 256'h0020000008800000000000000AA00A2000280A000A0808000A2020A020000AA0;
defparam prom_inst_0.INIT_RAM_3C = 256'h0AA02AA82AA8200020000AA820082AA80A2000082008028008200A202AA002A0;
defparam prom_inst_0.INIT_RAM_3D = 256'hC00000000000000020082008000820080AA802A80AA800080A0020A00AA000A0;
defparam prom_inst_0.INIT_RAM_3E = 256'h00000000000000000000000000000000000000000000000000000A0000002020;
defparam prom_inst_0.INIT_RAM_3F = 256'h2558000000000000200800000000000000000000000000000000000080000000;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[29:0],dout[3:2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 2;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'hF7CDCD13B007771D97A4E3DAFAEFAD92A2C234BCDB03039997EF3CD0F271F3EF;
defparam prom_inst_1.INIT_RAM_01 = 256'h093DBFCCFFB84BDBFD0B01E2FFDCBA3FCED2FC2F8D32BAEBBC307FD33A4E5370;
defparam prom_inst_1.INIT_RAM_02 = 256'h33BBB0EF2CF81C1FF22F2FFC71F2F364B487E7ECDBE1834FB55301EA380E6C1F;
defparam prom_inst_1.INIT_RAM_03 = 256'hD916FEBE0ADBF836BC032393BBFEF2E3FCCA08FFCAF8F4DCBC9BC17F8BCBF0F0;
defparam prom_inst_1.INIT_RAM_04 = 256'hEC701EE873EB454FE73EE25C6EAFC32BB95596AC243B55418D8C78C66477734C;
defparam prom_inst_1.INIT_RAM_05 = 256'h08027F73F52FCFC1C7E071D4B1E5B5965669B77568FB870E5722F7AFE3FCB0DA;
defparam prom_inst_1.INIT_RAM_06 = 256'h0F1377DC78000030003308383E435F8718CA343EEEFCDE3FBE36B7B08751E878;
defparam prom_inst_1.INIT_RAM_07 = 256'h3A38814400D050001C40440040040D7D48343EC24E020014840347BF354BDBF4;
defparam prom_inst_1.INIT_RAM_08 = 256'h8FC5E3EFE83EFE80D05E3EFE80C0FBFA30360D0501440DB924DFBFA33EFE8D58;
defparam prom_inst_1.INIT_RAM_09 = 256'hD1ECA2287FEE796F89D92D6C9E05286F64A1E2083100340711FB7C175B7A4501;
defparam prom_inst_1.INIT_RAM_0A = 256'h82008828400C04CB857E36E54539B87FA0361ECBE2FED2D8C703EBC1EB1527D4;
defparam prom_inst_1.INIT_RAM_0B = 256'h6E9371078B6D421E6E088CE0C0D124E9F87C04DC4E6E5D55623ECE36C6E1FF87;
defparam prom_inst_1.INIT_RAM_0C = 256'h94E9453615534231304043DC3C0CFEE6E1E348416364E9127D3CE000005573EF;
defparam prom_inst_1.INIT_RAM_0D = 256'hD1E19D0EB4BC86FA08718FA9FE8D92FC1C8FCF87A3D0D7DA345C4FB04F0D3BE4;
defparam prom_inst_1.INIT_RAM_0E = 256'hE7512E4860A6E0E04FAAB76A4DB064FB84A6A867347D4C498D12F2F7168BC83F;
defparam prom_inst_1.INIT_RAM_0F = 256'h355D50621B878B643F6CAD0B41778FD44D5550A9256AA7FFDDD8F9C5A276A243;
defparam prom_inst_1.INIT_RAM_10 = 256'h1CFDEBAE8F431368813C6D412B987F0ADAFCC2B58AD023A5AE2DADB0374CB254;
defparam prom_inst_1.INIT_RAM_11 = 256'hE9BE1A13204D9F92D6493BCEE89CAAD7D78FF4BA8F10783C1B5783AF22CAF7AB;
defparam prom_inst_1.INIT_RAM_12 = 256'hABBAEB000AA8AE6FC47BAFEA22290EF40EAABCAE2AD13B9316C68C850AC50BB7;
defparam prom_inst_1.INIT_RAM_13 = 256'hBD5BCAF838503BCB0FEB9CB422A2F35A82FA9A240A38E133CE8A7BC3483DB32A;
defparam prom_inst_1.INIT_RAM_14 = 256'hA38BAF361BC6F30174AD85392EAD8E3DAF8E82272FA9C4132BE0094A00A7AAF8;
defparam prom_inst_1.INIT_RAM_15 = 256'hAD8B9393280E351923B4933357B400001D82D4BE4D2CD8918034A04B8DBCEB14;
defparam prom_inst_1.INIT_RAM_16 = 256'h816F2FE68464B2344236B07F8C1401A3C256F9817BAA276EF8C7238A3C04EDBF;
defparam prom_inst_1.INIT_RAM_17 = 256'h4EE6E6DABA6080AC4F97BA03C9A8D7EFA0009D7AA0D8A00C8A34234236C4D558;
defparam prom_inst_1.INIT_RAM_18 = 256'h2C1221A12002A117BAD576A01A18BAFE9E1522BF59C080468AEB6AF9CA13E23B;
defparam prom_inst_1.INIT_RAM_19 = 256'hD43DADD1C9F9B453ACF80E3EBB68BB63FBEFE23A3AFA0C5021EB33ACCEFBA388;
defparam prom_inst_1.INIT_RAM_1A = 256'h28D8936884140DCE276F07C3487B53B32366E763F8C71BBBB8FC724E4E37EDAE;
defparam prom_inst_1.INIT_RAM_1B = 256'h6850DFA938C484E24256CE562DE77FD60A28FF658E7367B811A84A00539ACCB3;
defparam prom_inst_1.INIT_RAM_1C = 256'h8891BABB8BF797C5732F1F051E3DF077804FFBC3E73DE3689928461FD1E0004E;
defparam prom_inst_1.INIT_RAM_1D = 256'h0025EEFB8028A6B3FFA8D3BBA0CBF71EA7A4088C71C23D3FFE70D348E5F7E222;
defparam prom_inst_1.INIT_RAM_1E = 256'hF7C1A5FB14620DF6647F326E7237D6F6BB0EB8A30C74423B653E084FC121D8FB;
defparam prom_inst_1.INIT_RAM_1F = 256'hB4F81C02AAAAE950E60C4809C4764C785358A13F9C846BB891E3EAA9C76816CB;
defparam prom_inst_1.INIT_RAM_20 = 256'h1E27F38CAFFEBA8943FEC620BEE7B598328A801E0FEA13301311469FA90E1380;
defparam prom_inst_1.INIT_RAM_21 = 256'h0E6683C323FC0A88B3AFC2FD506AEC9B802812A80F144E639B43ECFA4FBDEE92;
defparam prom_inst_1.INIT_RAM_22 = 256'h6228890AA1A9397B2C8DD2A72A9A3604F7D020AA4EAAABBAEEABA4218D8DBB6A;
defparam prom_inst_1.INIT_RAM_23 = 256'h909638DA6BAC8E32AEA22892DE286ED6683983E0DE880001D9898698641F1686;
defparam prom_inst_1.INIT_RAM_24 = 256'h16AAA697078FE2A9606609ACA8EB10770AED14B30993020C8C50E73082A2828C;
defparam prom_inst_1.INIT_RAM_25 = 256'h9999C59999995A0C8C1DE00B800002088AEEAC9A608218593FD1E1E25C6F6962;
defparam prom_inst_1.INIT_RAM_26 = 256'hEDBDFF14053B4E2D27DDD987C0519958550119D15D929D512219955D9D5DDD99;
defparam prom_inst_1.INIT_RAM_27 = 256'hB01668276203101C1C0DFD47498B88CBB4C3DB837114AD8B6E4113844DADE28B;
defparam prom_inst_1.INIT_RAM_28 = 256'hF518A719B6DA0D030C78040030F69002E588397EA688B1E11A2035FA687172C0;
defparam prom_inst_1.INIT_RAM_29 = 256'hBE6E40911356F8433AF2D5F47A1AFE02A3978EF8BB6BEE3FF98019B8FFC8FD69;
defparam prom_inst_1.INIT_RAM_2A = 256'h2CA6E086C608872358DC8F74621F58F069A08E49BB926E669BA11351135B366D;
defparam prom_inst_1.INIT_RAM_2B = 256'h6F2F68DF3118DC67EBA8C101CEDE278D8C880C882376548D6391C651348D43A0;
defparam prom_inst_1.INIT_RAM_2C = 256'h746E23E2228DC5C8C700174DCBC3DEA3D37A17334FDC9E100BC1BCBF3813C13F;
defparam prom_inst_1.INIT_RAM_2D = 256'h24DE3B89BD0E746006D6483011AA1FA000022A44E8101403A228B1A82A76EA10;
defparam prom_inst_1.INIT_RAM_2E = 256'h40CFDD8AFC5C5A0CE34999CC104001901360084FF1009FB1E0B913E8397459E1;
defparam prom_inst_1.INIT_RAM_2F = 256'hC4030901123E3C7A433A6B0FCC86ECBD50C42C2402BA810284102330707237EB;
defparam prom_inst_1.INIT_RAM_30 = 256'hFFFFFFFFFA0411080149500E303A80EB172810EB700CEF86D9506853EBAD7030;
defparam prom_inst_1.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3A = 256'h02402800030028002BA01B9000001AA4000826201490BBB81D74001400000000;
defparam prom_inst_1.INIT_RAM_3B = 256'h224C09800CC0189000000000330C30CC024C30CC30CC2EA830CC330C3AA8309C;
defparam prom_inst_1.INIT_RAM_3C = 256'h300C060000903000062430003AAC00C0330C00CC30CC2418300C30CC030C336C;
defparam prom_inst_1.INIT_RAM_3D = 256'hC0000060000018003AAC309C00900690180024003000000C30CC070C380C030C;
defparam prom_inst_1.INIT_RAM_3E = 256'h256015601560300018209544200015809D70008C326035D4303030C03760308C;
defparam prom_inst_1.INIT_RAM_3F = 256'hC823002400C02AA83A2C30B09D50189025500A5025503020262000305D700960;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[29:0],dout[5:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 2;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'hD442423B30A09C2C532B0ADBD3C32F550FA2CC342C6C6C1DD7510426B5781070;
defparam prom_inst_2.INIT_RAM_01 = 256'hB2CF35298050C3F35263B242D522BE808100D35D0883DB426200F21032B09045;
defparam prom_inst_2.INIT_RAM_02 = 256'h9B321E11094290BC81B30C8CF61A7E2B3AE9E96AF35B9B30CFF0227CB008C79C;
defparam prom_inst_2.INIT_RAM_03 = 256'h31EDDD743BFAD6C83EA9642C00D51F2B5668820706CB01B6669562F5ACC35A7A;
defparam prom_inst_2.INIT_RAM_04 = 256'hF002034EEA73182873A332AB2CCD2433CC00C3D5B73C0020CD8058147754D0B4;
defparam prom_inst_2.INIT_RAM_05 = 256'h92204F34F0A1C80A20A0B4C28802E08A03AE99D8B5B13228036CD4503A12FCC8;
defparam prom_inst_2.INIT_RAM_06 = 256'h07A94A52FC2B2C0800290C233F2E2CC23EA7233FE984242D300B6404640904E8;
defparam prom_inst_2.INIT_RAM_07 = 256'h370A80A2020A20020722A2C02C0088B2CC233FCA228AC02CC0FD22610AC60ADA;
defparam prom_inst_2.INIT_RAM_08 = 256'hB80B32A1FC2A1FC084B32A1FE028A87FC82300A200A2E9783A0A87F02A1FC8B4;
defparam prom_inst_2.INIT_RAM_09 = 256'h0043857683233C378504113CC785231663F803048CC012C1C2A8FCC38E4E080F;
defparam prom_inst_2.INIT_RAM_0A = 256'hB0514185C04C0D2A640DB2992126DA80D05E80C342D70AE2CCEB40C320087526;
defparam prom_inst_2.INIT_RAM_0B = 256'hCAACB2490BB292CCC793AEFAD6DB6B3A06800A6C822E822666E26A398BAA00E0;
defparam prom_inst_2.INIT_RAM_0C = 256'h0A0682892B2892C007C0CC53118006CC7A0B9482FA2B0752B72A3C8C00C7CAA1;
defparam prom_inst_2.INIT_RAM_0D = 256'h44459CC466AD4AB137C8CDF919B170D6F2E3E44CAE68A06A8E50064AB3CDE0DA;
defparam prom_inst_2.INIT_RAM_0E = 256'h039B0F44C2CC79408BC7E3B2B152C2BDE04BFD0A8352603691B0CADB230EF0DC;
defparam prom_inst_2.INIT_RAM_0F = 256'h8986A4C2F1E90BD8ADB1AE6B8BB9182EB0000000000000CCC4888AC8C2771C27;
defparam prom_inst_2.INIT_RAM_10 = 256'hA2B62BA2B9A201AAA22FB1A1A8884F8AEA159689440068B9A0B6A243100196A8;
defparam prom_inst_2.INIT_RAM_11 = 256'h4B4CACAC24B0A4F0EDB1E03821AF2AE869181C33EFA49296ACA52925A50ADB68;
defparam prom_inst_2.INIT_RAM_12 = 256'h68A2E8AA9BE2A223E2FA2F48C4B638195182B5C12709E04B3EEFAD697EF1AEBB;
defparam prom_inst_2.INIT_RAM_13 = 256'hA228DAD23EA09569E3AB2EB2C6CAB9A6AADA82C2A81B288B2C2C2395AB0668A1;
defparam prom_inst_2.INIT_RAM_14 = 256'h690B239978363904E5AEB2C30FAE91ACADB2082CA80B01A02B41B2ACD12C1E0A;
defparam prom_inst_2.INIT_RAM_15 = 256'h85782C19A1872A8BF54DACD0E61ABBBBB68E0C38B30D0AE8C06A9BABA7832BA9;
defparam prom_inst_2.INIT_RAM_16 = 256'hF8CDC929412C31280B2A8AE48D3D5BFBE60549A9496E0BB82637773EBE006334;
defparam prom_inst_2.INIT_RAM_17 = 256'hAE66226896EFB2B804949601282B3927600880BA8B93E938BE80C2AACBAE51E3;
defparam prom_inst_2.INIT_RAM_18 = 256'h38B2C36BB3B803949608556A2B2EBAB6B2A8A983A88B0203061C0D8930AC42C1;
defparam prom_inst_2.INIT_RAM_19 = 256'h20ACAEC2C8E6C02A3A1C2BA46486E4AAEC2BA026E6B8836058CF7B5DCDE43BBB;
defparam prom_inst_2.INIT_RAM_1A = 256'h8CA7CECBE0C08B3CFAC16F8C34CC2268FACBAC059EC0D643F7E0223BB924B039;
defparam prom_inst_2.INIT_RAM_1B = 256'h9C029BE1FC0F0F8CF20DA3819BAC21549C31AC26CB8A2BE23B8EDBB8E018E5B8;
defparam prom_inst_2.INIT_RAM_1C = 256'h52017C6C9602F1A06077182CB6B5DBA4E0BA0DB5B60DFA55504B2B4B0AF020B9;
defparam prom_inst_2.INIT_RAM_1D = 256'hAD118360C095133FE470936CB886F3FCC5B98803FFD480AB28196A9E2E306944;
defparam prom_inst_2.INIT_RAM_1E = 256'hC28EC4E005937DB0BD60B2B127662BF33DA62672FFF0F4F32B0EC0336B5FF33D;
defparam prom_inst_2.INIT_RAM_1F = 256'h54A4C1351144841EC8B664956656220EC8E0F70BB0000B3223C716694A5406C6;
defparam prom_inst_2.INIT_RAM_20 = 256'h2DAE4336998E296AEE4B1E33C9224967461ABBB4802288BA99A9ADB885251101;
defparam prom_inst_2.INIT_RAM_21 = 256'hC25970B44600BCEB88BB0AB19AD2CA780D34D4382343495E3530B42D42DCB6B9;
defparam prom_inst_2.INIT_RAM_22 = 256'hD4451067189BAF2C988EDDDD9C4CBAF377E2386695144511445653586A6AEC9E;
defparam prom_inst_2.INIT_RAM_23 = 256'hBDCD65A196535967699445154A9A9B25970BF0AD0065BBBB51C569B452C0D596;
defparam prom_inst_2.INIT_RAM_24 = 256'h32CCC292E7183530245310C0B0299926F5EFBEA32BA3A99D6CCCCBF1E14D3556;
defparam prom_inst_2.INIT_RAM_25 = 256'hFFFFB7FFFFFFB77B33BF0324330C307BBA440F88158CAD3BAB12ED06ED8F08B6;
defparam prom_inst_2.INIT_RAM_26 = 256'h16EC00A73AB59996FF33B7363B737F3F33B3337FBBB73B37B3F7BFF7BB3F77FF;
defparam prom_inst_2.INIT_RAM_27 = 256'h005CB542198E064D4E2EC00B2678A3B819B06619002456F1896E994B5845F137;
defparam prom_inst_2.INIT_RAM_28 = 256'h772E2B0781C32B00E30C22C80F40B5B6102B0B06A8670F1CA68B0C1A40000DF7;
defparam prom_inst_2.INIT_RAM_29 = 256'h7DE0C8FBBB08280C1C8EC0F7775381AF2C0AA528141E50601920578180BEB24B;
defparam prom_inst_2.INIT_RAM_2A = 256'h4A352D75F232EFAC1B3370C24E7CB33241C5595B8966E29DB88BB9DBB38AA1E0;
defparam prom_inst_2.INIT_RAM_2B = 256'hB30CEB956B1B3639602B1F0323905BD6B8BE38BE2CC01AB06C313F7F1FEBB16A;
defparam prom_inst_2.INIT_RAM_2C = 256'hDA9A2CA12FB3C52B1C301842595750AC069654A843E5A5B0256ACC359022F88D;
defparam prom_inst_2.INIT_RAM_2D = 256'h32938FF5F9FAAE8E8B69D08C2CBBFE320C83CF0F8E00A2C219C66A554557518A;
defparam prom_inst_2.INIT_RAM_2E = 256'h12B76B06DEB794AB653651908BF220DFF2F080C00FC0FA83F20C3F8E23234C0C;
defparam prom_inst_2.INIT_RAM_2F = 256'h33CA340BC1A33F4321E325B81AE6B2164233F8D08AE34308C03CACCC8B23AF8C;
defparam prom_inst_2.INIT_RAM_30 = 256'hFFFFFFFFF3808320F30C83CB93E34A8CE0A48F8C0EBE597EF382E6F1D7D24742;
defparam prom_inst_2.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3A = 256'h2400140003004000030013102558000000103264092833B02EB8002811540000;
defparam prom_inst_2.INIT_RAM_3B = 256'h000C10100CC0010094101040330C30CC140C30CC30CC0C90300C330C3024390C;
defparam prom_inst_2.INIT_RAM_3C = 256'h300C00600060300000C03000300C00C0300C00CC30CC300C300C30CC030C314C;
defparam prom_inst_2.INIT_RAM_3D = 256'hC0001574355C01800000390C15800960240018003000155C30CC030C310C030C;
defparam prom_inst_2.INIT_RAM_3E = 256'h30300030156005542BE8600035C400C0CC301550333030C01A903AE833303AE4;
defparam prom_inst_2.INIT_RAM_3F = 256'hC6930024351C000000C03930CC00098025401A003000057433302A900C300C30;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[29:0],dout[7:6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 2;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'hCB3E2FC3EC07CFCC3000C0C0FCF3CF30C93CF4F3CFC7CFF7702CF2F0B000CF1C;
defparam prom_inst_3.INIT_RAM_01 = 256'h2C38F0CB2C0B4FCF0F0F2F2CF3F03C1C73E3D8819D0094673CF031C3000F830C;
defparam prom_inst_3.INIT_RAM_02 = 256'hC2DED43D9C303C0C302E3C3C32D44704FC0D0D404F510000436007401C0FB50B;
defparam prom_inst_3.INIT_RAM_03 = 256'hFFFF3FF2F0F0FCFF740143C33CF1D40FD4533C73C0F2D5C5750140350BCF5343;
defparam prom_inst_3.INIT_RAM_04 = 256'hD50081B46AA05C07A01D5032040D830350000106103500004D0CC0CFDF4BCFB2;
defparam prom_inst_3.INIT_RAM_05 = 256'h1E075D70C12D5C73C30CF044B0F350BE016F88093E8D430703E0CBC011D860C0;
defparam prom_inst_3.INIT_RAM_06 = 256'hF51CBD2D30EC30CC0CF3F030B433C70F82E030B40CF2F2CFF303CFD743D0CF48;
defparam prom_inst_3.INIT_RAM_07 = 256'hB00330F3330F3CCC3023F3033030CF1C7030B40C30CC0CC700002F3CBC73C0F0;
defparam prom_inst_3.INIT_RAM_08 = 256'h0C72C30D4030D400F32C30D4333CC3500CFC30F330F33C00CF3C3500F0D40F1F;
defparam prom_inst_3.INIT_RAM_09 = 256'h70CF3F1CF40085953F43F60821435E06D090FC30800CC20C03C3F00FC0F00C00;
defparam prom_inst_3.INIT_RAM_0A = 256'h2DCF00C0C0A3FC0A0010008FD1735BC040100F4F2CF1C0FCC7C32CC1F102D3C8;
defparam prom_inst_3.INIT_RAM_0B = 256'h5C032C3CB33F0CB7B4330C70C07F00F0300C0CCFCEEAFAA660C400D5CD6F4043;
defparam prom_inst_3.INIT_RAM_0C = 256'hF0D32C33F0C30CB003C0C3400C00B07B4033C43F0B00C1309572C08206000B0D;
defparam prom_inst_3.INIT_RAM_0D = 256'hF02C0CC2EC2C003300B03D02C32C33D42CC34C073B51E053001C0CB00C1D0B0C;
defparam prom_inst_3.INIT_RAM_0E = 256'h4CC13DF3B07F432DCB4034D00F8070F50C382743103C84331C13C0F3FEC3EC3D;
defparam prom_inst_3.INIT_RAM_0F = 256'h13DFC3F0ED0CB3CC0F3C0F03C33CB2F00C0000003FFFFF33373330FFF03C0F03;
defparam prom_inst_3.INIT_RAM_10 = 256'hF03F032CED47014F072F3FC00B010D10F2D5FCBB32F00C232C2F2F30CBCC14FC;
defparam prom_inst_3.INIT_RAM_11 = 256'h501FF403470C2423FCEC0B02FC0FC0FD3CB2FCFF0D03D0D4CFFD0D053CC0FE0B;
defparam prom_inst_3.INIT_RAM_12 = 256'h0B3CCB00026C2C0345D3CD4373F302FFF0F03FFCF2FC0B02BC8F0C0FC038081D;
defparam prom_inst_3.INIT_RAM_13 = 256'h3FF3D0F0F7F011430F43F03074703FC3D0FF007401F2F11007476CBD4CF5701F;
defparam prom_inst_3.INIT_RAM_14 = 256'h14B30FFD73F0FF03ED0F3C3E3F0F1F0C0F2F50CFCFC3C0F303D41F478F0F00FF;
defparam prom_inst_3.INIT_RAM_15 = 256'h30CBC3D13FCD7BC09CBC03CBFED411111532F8FB0E3F50E0007B0FC35F3F03FC;
defparam prom_inst_3.INIT_RAM_16 = 256'h413D5D4C0004F4780C3CFCE530BC03C3404C53C07144F3C2F003030C340044F5;
defparam prom_inst_3.INIT_RAM_17 = 256'h44444453144D1CECF50714014333F94C3C0F3FD03EFE7FEC27D407BCFEC05FFE;
defparam prom_inst_3.INIT_RAM_18 = 256'hEF0070151D100D07145FC30005F83C3F3D73C33F3C01C0C3F3CBC0F2EC032CBD;
defparam prom_inst_3.INIT_RAM_19 = 256'hF00C0FCDC1F3032F00F0ECB2C3C003C0C3030D732DCC0CF003F7C7DF1F03F011;
defparam prom_inst_3.INIT_RAM_1A = 256'h30F303C33000FF03CB0D8C00307023C3CBF8CB5590C13C3C3CC7700B8BCF0FC0;
defparam prom_inst_3.INIT_RAM_1B = 256'hF0FEF00F000000FF300F2C0A0CCB6587F55E877F0C0B093F01A4691030DA4691;
defparam prom_inst_3.INIT_RAM_1C = 256'hCCDBDFCBE0775984CF03B3F6160818CF330C758984F74F4FF0420901D243330F;
defparam prom_inst_3.INIT_RAM_1D = 256'h8CFD2D4B400CF035CFFC28CBCCD1B04C0D8C01C134C0001F1C1862CC04906333;
defparam prom_inst_3.INIT_RAM_1E = 256'h172E5D0701C703039C3C109047A3E0F035867FC35D3030030934D01763C4D175;
defparam prom_inst_3.INIT_RAM_1F = 256'hD42F0FF0CF333DC0FBF44FFF44D744D451FF71310500F3DCE07D440141C30C00;
defparam prom_inst_3.INIT_RAM_20 = 256'hB700F003F8677F177CF2EF5092F4BFFCBCF011180CB3D110113308C7FC03CCC0;
defparam prom_inst_3.INIT_RAM_21 = 256'h3FFFCF8BFCB4243CBD91DF1FF08CF8CFFC000300050C7B72CC0314C74C51D013;
defparam prom_inst_3.INIT_RAM_22 = 256'h333CCC0DF001010FB822437537C0090700209FFFC0F33CCF33F7C000DFDE4BD3;
defparam prom_inst_3.INIT_RAM_23 = 256'h33C37DE0B7C0DF70DF333CC0C975F2FFFCFF0FB2CFFFD1110C7FCC0E300C0CCC;
defparam prom_inst_3.INIT_RAM_24 = 256'h003334F7EDF2F0CD0810A0F01C0112CC000C10280228002D0002F90E7F3CF5D7;
defparam prom_inst_3.INIT_RAM_25 = 256'h0000000000000048C080826C700923D113333C0E1418261121FE72FF6C3C40F0;
defparam prom_inst_3.INIT_RAM_26 = 256'h03570074BB1D5FF512C0004848088C04C88C0C08884848C0C40C884C4448C800;
defparam prom_inst_3.INIT_RAM_27 = 256'hF03FB0327FFB00807403443DFFCB5ECBD5CF57FC303F353D5FF11100C4C5F303;
defparam prom_inst_3.INIT_RAM_28 = 256'h02B4090CF0CC3C301CF0F338C077F01340FCFC353FFCF3F33D7CF0D4F0181C3C;
defparam prom_inst_3.INIT_RAM_29 = 256'h333F3F62217CC30195C2EA0030B02C090FFC02C30B072FCB60C03CFF2D271FF1;
defparam prom_inst_3.INIT_RAM_2A = 256'h0C08083030E079CFF3F003C07FC3F000737C08FCFF2F3FC3CFFD104110C2203C;
defparam prom_inst_3.INIT_RAM_2B = 256'h3E3C0EF57F33FBDD43F2CF03003FCFC52C27EC27CBD4FF3FCFC333FC3F2FBF0C;
defparam prom_inst_3.INIT_RAM_2C = 256'h14F0CF0C093CB0F2CC000F0F50B32FCB5794C3CF0F353530214CFCF50B72FC0F;
defparam prom_inst_3.INIT_RAM_2D = 256'h003CFD369CA32CF195950880C008C3C200CC3000F30CC30FFFFCF2003C617F03;
defparam prom_inst_3.INIT_RAM_2E = 256'h2875ACD3DEE8AF95A9C6D088800220C4C300800FDC000C38423000F23D7080C2;
defparam prom_inst_3.INIT_RAM_2F = 256'h000B000800B0B4BC003C313F2C93CA0722000C00C83C000B00C08000081B30F0;
defparam prom_inst_3.INIT_RAM_30 = 256'hFFFFFFFFFC80802000F0000C803C08F0008080F00A79FD1382F5BE42E61B4222;
defparam prom_inst_3.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_3A = 256'h0000000000000000000000000000000000000400101400000410000000000000;
defparam prom_inst_3.INIT_RAM_3B = 256'h0010000000000000000000000050051000040550045405000410141000000550;
defparam prom_inst_3.INIT_RAM_3C = 256'h0550155415541554155405000000155405501554155415540550155415500550;
defparam prom_inst_3.INIT_RAM_3D = 256'hC0000040100400100000100400181004055401540554000C0410155405501554;
defparam prom_inst_3.INIT_RAM_3E = 256'h0540155015500000000000000000155401400000054005000000000004001040;
defparam prom_inst_3.INIT_RAM_3F = 256'h1AA4000010040000000010100150101005500050055000001040000001405550;

endmodule //Gowin_pROM_1
