//Copyright (C)2014-2025 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.11.03 Education
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9
//Device Version: C
//Created Time: Sun Sep 21 11:06:49 2025

module Gowin_pROM_test (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [12:0] ad;

wire [29:0] prom_inst_0_dout_w;
wire [29:0] prom_inst_1_dout_w;
wire [29:0] prom_inst_2_dout_w;
wire [29:0] prom_inst_3_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[29:0],dout[1:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 2;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h92ED8B62B8A62B8A18170F0DE0C9D3B1A7DE7BFFFFFD1341291554140037AFA7;
defparam prom_inst_0.INIT_RAM_01 = 256'h1B302CE0E00552E0A0C886E2B105C155C115013D1D75B65B702619AAECBB2E9B;
defparam prom_inst_0.INIT_RAM_02 = 256'hC121F742054854C490555096328957245F7FE32212550B0245480E8454B02056;
defparam prom_inst_0.INIT_RAM_03 = 256'hEF9EEAF9545754E4FCB279E4400E5652FB7750515CBA2BFC3954957854846DD0;
defparam prom_inst_0.INIT_RAM_04 = 256'h02ABFFFEA801561520B6BEB3BF292E5641061F408A45405E1425505520922BE7;
defparam prom_inst_0.INIT_RAM_05 = 256'h315C1C156545F4529125730715DC2CB9D81C1D57D711169C450AD91A54015554;
defparam prom_inst_0.INIT_RAM_06 = 256'hE14A56143CA30BF26381510FB3FBFB2E284FFC1DFEBE14124E0454509544BBF7;
defparam prom_inst_0.INIT_RAM_07 = 256'h4BEE9512EB8EB14A060456F85095715051214A55C541C2E8E24377C3CBC3CB81;
defparam prom_inst_0.INIT_RAM_08 = 256'h957B2EF7093BE0D1A09DED2481BE075624823A02C0AC24A0944E054263E8BBBA;
defparam prom_inst_0.INIT_RAM_09 = 256'h46AC6646042AA298281CEA4E85079545E5515C7DB900AFB5C702BED6291514A0;
defparam prom_inst_0.INIT_RAM_0A = 256'h7FAF619F2FD6C1C1067F6F619F2FDEC1C1067FEF53CF41150410954155488245;
defparam prom_inst_0.INIT_RAM_0B = 256'h5019FD0619E2FDF070419FFF7070719C28B07DC1C1467E2C1F619F2FDAC1C106;
defparam prom_inst_0.INIT_RAM_0C = 256'h410410550454104A55679B99A6265545095612A4E56507C57549914A5567127F;
defparam prom_inst_0.INIT_RAM_0D = 256'hD68356C2356982B6A0456F8509544A45654141C85510410507F8A041052FD868;
defparam prom_inst_0.INIT_RAM_0E = 256'hA041BE44954E428C0757D2C5BE7C1D7EB9B1FF3B4F2E0BC773B407FFEB2FE601;
defparam prom_inst_0.INIT_RAM_0F = 256'hC0757075F3E80FF2C4C7F24CFA4C4D3F4FE3FCFFE9CFB106C9ECA3B17876FB7D;
defparam prom_inst_0.INIT_RAM_10 = 256'h46F4ACA0456B6CB2DBAD45DD0B1BE142556FBCDB103FCB131FC9CFB0F0FD3F8C;
defparam prom_inst_0.INIT_RAM_11 = 256'hEC460ABD444B5046FC3BED7F43BAF733A6F4BB6BD041BEC554E42E027DAF61D0;
defparam prom_inst_0.INIT_RAM_12 = 256'h3F51D619CB5E503BEFAF457F523EA507E2FA2E7620EEF5152D5721562C612C1B;
defparam prom_inst_0.INIT_RAM_13 = 256'hE3D6FFCB77743E8B440FF98AF64726F8E3F2173FD85E1DC8A3590763F3191D70;
defparam prom_inst_0.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000001F6B95E627FEBFA0BFFC59;
defparam prom_inst_0.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_20 = 256'h060A0D51F6355C6271E0D0537E51634C22539C4393CE470A7602F6512EBAB422;
defparam prom_inst_0.INIT_RAM_21 = 256'h7C2C134160A04D034824134273C2013409F0B04D092E0A04D02797090D5940D0;
defparam prom_inst_0.INIT_RAM_22 = 256'h4A0606460045343D3782C1343BC60904D0BB82013424980824134107DC201343;
defparam prom_inst_0.INIT_RAM_23 = 256'hD031110213105974040C840C841653409E5C58D30B9D20039762539CC5E99F09;
defparam prom_inst_0.INIT_RAM_24 = 256'hCF635D725330D68C5CF63C55D7100D0FB95D23122230230597440C80C80C4165;
defparam prom_inst_0.INIT_RAM_25 = 256'h09F06BCB132F70435012E079139A60D0D019407AC43424B816B044C35A309331;
defparam prom_inst_0.INIT_RAM_26 = 256'hDE3A5BC404F01C5C841B39F60401634CD0701341249808407F3424980890C434;
defparam prom_inst_0.INIT_RAM_27 = 256'h04036BF410467DD896136BC04CD67C100C4C58D3341309260210DAF0E31479A7;
defparam prom_inst_0.INIT_RAM_28 = 256'hD2643698D09CF216E2498100CCC35A3D838D0D030A4610492604036BC410509F;
defparam prom_inst_0.INIT_RAM_29 = 256'h4027305C040F61841C34F3414DCBBB9451365F056F976F96DBD2756F19BD49BF;
defparam prom_inst_0.INIT_RAM_2A = 256'hD8446441976305C440F618490D16A93939393939390162718C11161602411113;
defparam prom_inst_0.INIT_RAM_2B = 256'h2540C350DAF25841C3453414DC41F7A3CD034A8CE45C4024C35A3D8BAA805865;
defparam prom_inst_0.INIT_RAM_2C = 256'h0402763E59B09140BDC79475305CC40F60B62F60914393D801B47C1100729849;
defparam prom_inst_0.INIT_RAM_2D = 256'h7C110072D972103D82A1072540C250DAF258490D16493804BD8DC6C107D30911;
defparam prom_inst_0.INIT_RAM_2E = 256'h994E45C403330D68F616AA009A50477D4F1001D278D1B0409312D650E7D801B4;
defparam prom_inst_0.INIT_RAM_2F = 256'h1980010D201980011DA10DA11D780101C10D780101C11D4903662424EF343D37;
defparam prom_inst_0.INIT_RAM_30 = 256'h309E25330D68C5CF62FD37840343E6F151382F00C10D382F00C11DA101A11120;
defparam prom_inst_0.INIT_RAM_31 = 256'h0D68C5CF61E92CE7BC95B54B30341634CD033416230D04024CC17193D8F34162;
defparam prom_inst_0.INIT_RAM_32 = 256'h06492807531601924001D7AD1F16C51166D51058D058D3340C45834A30D01463;
defparam prom_inst_0.INIT_RAM_33 = 256'h17193D833437F9C340518C35A3173D8BB51836BC4067A553BA4E7D8124E34C58;
defparam prom_inst_0.INIT_RAM_34 = 256'hC458D3643930DCB44C4645E84439F0E1009CC61070D14D05373BC6A0D04024CC;
defparam prom_inst_0.INIT_RAM_35 = 256'h8ECB44C7A11065D8C6124345AA4E4E4E4E4E4E40589C630445970107D80ECB44;
defparam prom_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000E45C4024C35A3D85AA805865D8445971103D;
defparam prom_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3A = 256'h002000000200000002000200000000000000220028082A200820000000000000;
defparam prom_inst_0.INIT_RAM_3B = 256'h0020000008800000000000000AA00A2000280A000A0808000A2020A020000AA0;
defparam prom_inst_0.INIT_RAM_3C = 256'h0AA02AA82AA8200020000AA820082AA80A2000082008028008200A202AA002A0;
defparam prom_inst_0.INIT_RAM_3D = 256'hC00000000000000020082008000820080AA802A80AA800080A0020A00AA000A0;
defparam prom_inst_0.INIT_RAM_3E = 256'h00000000000000000000000000000000000000000000000000000A0000002020;
defparam prom_inst_0.INIT_RAM_3F = 256'h2558000000000000200800000000000000000000000000000000000080000000;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[29:0],dout[3:2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 2;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'hD6309C6F19CEF19FBC7BBA8BE3A76B7BF3CF86FFFFFC91070833EF0C001FF1DC;
defparam prom_inst_1.INIT_RAM_01 = 256'hBD9A3438368CB33C362E4331901E4737802E801170C71CF1E9EFB9DA33ACA37A;
defparam prom_inst_1.INIT_RAM_02 = 256'h60B370D1028F0268682AA85204E6AB1C0B3F59199156AF9382CFA7282CD93C2E;
defparam prom_inst_1.INIT_RAM_03 = 256'hBBEFB7BE2FEEEA286DC331FCF40FB231C7EED0002054AFFDB70C71F70C78CC36;
defparam prom_inst_1.INIT_RAM_04 = 256'hA80154015555578B38F1DDD07F1E1C41C002AE8AA0C0E1EF2C63E84B3AEF1EFB;
defparam prom_inst_1.INIT_RAM_05 = 256'hE03828001D40F0B28F33DA1E03FF325ECC0478DFC93320C40B2B0CF73C02A802;
defparam prom_inst_1.INIT_RAM_06 = 256'h72CE3D81A1E167F1E1742308A3AA2293304E6B0B607394014F1C0CB38FA2A22E;
defparam prom_inst_1.INIT_RAM_07 = 256'h2C721535FCC4F0CF2B1C0F1CB18FA833CFB2C23EA0CF835079899DB045B044E0;
defparam prom_inst_1.INIT_RAM_08 = 256'hCF9C95F8863EF97371F00B6347C7842F63429F3B02706F61B87B1487C3C47ECB;
defparam prom_inst_1.INIT_RAM_09 = 256'h2BB6F7E741AEEBDC9C06BBE701634115C403682D7FEC79D06CB1EF4383032C6A;
defparam prom_inst_1.INIT_RAM_0A = 256'hD4BF1A3633C78780A8D47F1A3733CF8780A8D4FF362F07033C728FA30B5CE3DA;
defparam prom_inst_1.INIT_RAM_0B = 256'h39837CC1A3633CE1E02A353F21E00A3538403C878068D6100F1A3533CB8780A8;
defparam prom_inst_1.INIT_RAM_0C = 256'hC00003CF1C0CF1CE3E1F8F47E312CE0B38F4960C40DBC062E2E082CA3D1220DF;
defparam prom_inst_1.INIT_RAM_0D = 256'h5EE17F4C17A4F0D231C0F1CB08F660C0DBA302A40E3000010A00E0000211C02C;
defparam prom_inst_1.INIT_RAM_0E = 256'h91CFC74BCBCB23A461B40182C79878D37CF2BA0AD435A782E0AD313CFC3F9B8F;
defparam prom_inst_1.INIT_RAM_0F = 256'hA9EAA1E97B3C2961878AA18ECF747B9645A16C5B3EAA00330E7059E0B22D02C0;
defparam prom_inst_1.INIT_RAM_10 = 256'h9F303231C0E41041041A0C03460C72C23E31DE0600A5861E2A87BA106C581644;
defparam prom_inst_1.INIT_RAM_11 = 256'h70AF06E00AEE889F37075A1B3079820D938242E401CFC784B0B63343E09012B4;
defparam prom_inst_1.INIT_RAM_12 = 256'hB610B9A747EE3306666809F82C19A31E23A23A223C15E027B82E2273182B90FC;
defparam prom_inst_1.INIT_RAM_13 = 256'hC020AD8ECECC33CC986DB6CD438EA16C96214FB6CC872B6CD9ED82DB61A70BB8;
defparam prom_inst_1.INIT_RAM_14 = 256'h000000000000000000000000000000000000000000243B072415D257F153D80E;
defparam prom_inst_1.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_20 = 256'hF50C04F80413D58403C114D480F34440A08CE06432C793C88BBB644472021230;
defparam prom_inst_1.INIT_RAM_21 = 256'h3034345300D0D148343434507F0343451DC0C0D1414C0C0D1443260C04E72114;
defparam prom_inst_1.INIT_RAM_22 = 256'h8C48140400E345224B83434523570C0D140003034505E0283834515400383452;
defparam prom_inst_1.INIT_RAM_23 = 256'h40321210110213D0088444400084F4510C98D110283435C804408CE028C3C7CC;
defparam prom_inst_1.INIT_RAM_24 = 256'h004132601C348408E004123F26191147D3F40033010220213D04C8884440084F;
defparam prom_inst_1.INIT_RAM_25 = 256'h1DC22008007C40041C40D20301EF411429147201004505308841A4D210216800;
defparam prom_inst_1.INIT_RAM_26 = 256'h484F500648C3E49886771E04064F444029F4581405E02809904505E02A310045;
defparam prom_inst_1.INIT_RAM_27 = 256'h06447F0930F8011C6F547F0F902C5C1913A4D1100A7341780A011FC1F37E1EC1;
defparam prom_inst_1.INIT_RAM_28 = 256'h0CCD9811141FC4CCF05E0190D0D2100104D142934C5430F17806447F0C3D1C17;
defparam prom_inst_1.INIT_RAM_29 = 256'hA4743498064043945C4504535200013CD69CF7F6C0C8C0D4700753C053017302;
defparam prom_inst_1.INIT_RAM_2A = 256'h1011F111644349886404394E117FFA95403FEA9540FFE7410D047F5001840470;
defparam prom_inst_1.INIT_RAM_2B = 256'h0630D0B11FC33945C45F4535205500401148361079846474D2100100FE3FF959;
defparam prom_inst_1.INIT_RAM_2C = 256'h4647941FFDF41471F10430633498064040CF4C41C230301035F98C1049933D4E;
defparam prom_inst_1.INIT_RAM_2D = 256'h8C1049933E6219010335170630D0111FC3394E117FB13015310047D19E181C10;
defparam prom_inst_1.INIT_RAM_2E = 256'hA3C7984643434840043FF8FE3C100501CB193E777421F464D92FFF8C0C1035F9;
defparam prom_inst_1.INIT_RAM_2F = 256'h1240C804001240C834C804C834700101F804700101F834DC998872570045224B;
defparam prom_inst_1.INIT_RAM_30 = 256'h410C01C348408E0041224B864451F408F0703741F804703741F834C800C83000;
defparam prom_inst_1.INIT_RAM_31 = 256'h48408E0043314C7A34EE3DC72002344402944530C411464410D262C01004530C;
defparam prom_inst_1.INIT_RAM_32 = 256'hD45D1499F044351740267F3E43FE3857F8F7274408D1100A5178445841144443;
defparam prom_inst_1.INIT_RAM_33 = 256'h262C01044523210451100D2102380100C5C4443064594E303047811425F4C110;
defparam prom_inst_1.INIT_RAM_34 = 256'h0CD110C67C3444F910C46FC4111E7FD191D0DE517117D14D482357411464410D;
defparam prom_inst_1.INIT_RAM_35 = 256'h044F910F10445910DE53845FFEA5500FFAA5503FF9D043411FE6019C10344F91;
defparam prom_inst_1.INIT_RAM_36 = 256'h000000000000000000000000000079846474D210010FFE3FF9591011FE621901;
defparam prom_inst_1.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3A = 256'h02402800030028002BA01B9000001AA4000826201490BBB81D74001400000000;
defparam prom_inst_1.INIT_RAM_3B = 256'h224C09800CC0189000000000330C30CC024C30CC30CC2EA830CC330C3AA8309C;
defparam prom_inst_1.INIT_RAM_3C = 256'h300C060000903000062430003AAC00C0330C00CC30CC2418300C30CC030C336C;
defparam prom_inst_1.INIT_RAM_3D = 256'hC0000060000018003AAC309C00900690180024003000000C30CC070C380C030C;
defparam prom_inst_1.INIT_RAM_3E = 256'h256015601560300018209544200015809D70008C326035D4303030C03760308C;
defparam prom_inst_1.INIT_RAM_3F = 256'hC823002400C02AA83A2C30B09D50189025500A5025503020262000305D700960;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[29:0],dout[5:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 2;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'hC4330CC311C0712F8CC19EC27F0789AEF3DA3FFFFFFF618C48C23D2C000BF4DB;
defparam prom_inst_2.INIT_RAM_01 = 256'h8DA500B239E48B923D8C23B49030EF9982014010430C100134C732C0B01C0710;
defparam prom_inst_2.INIT_RAM_02 = 256'hD2FE715308EC60C0146AA88365C0AA243A002E36F9243E40E22CF7DE22C40220;
defparam prom_inst_2.INIT_RAM_03 = 256'h37C77F7CE42532F280D600CE000310900ACCF2422300CD544B23B20B23B38C54;
defparam prom_inst_2.INIT_RAM_04 = 256'h6F906F906F906F48B1C012C015ED14A3010A9778A013031D31220E48B3CFBDF1;
defparam prom_inst_2.INIT_RAM_05 = 256'hC4CEF0093181F8048C7216BE4C63750B1C2EFA67E10E20A4404B5CCF23906F90;
defparam prom_inst_2.INIT_RAM_06 = 256'h3012236274F639E8C8BA28DDFDD444098FEC37CC7493C820E73130C4885AC444;
defparam prom_inst_2.INIT_RAM_07 = 256'h5D32E3A82DD0D2A7A331334CC5883CC30CF01620F30C6312B0AEC336D336D012;
defparam prom_inst_2.INIT_RAM_08 = 256'hC83D322FAA5DF0BB744100404CD3E62340520EF3AF3B112C4EFB46F10B0E9DD3;
defparam prom_inst_2.INIT_RAM_09 = 256'h23023023018C18C28C0A30A30104AC1E408CBD44336EF7C25CBBDB1A804C3163;
defparam prom_inst_2.INIT_RAM_0A = 256'hAEBFBC2BBBE7EF82F0AE7FBC29BBEFEF82F0AEFF821F0C4C30C58839C8C6C700;
defparam prom_inst_2.INIT_RAM_0B = 256'h8BD2BE4FC2BBBEBBE0BC2BAFBBE0BC2AB4607EEF82F0AD181FBC29BBEBEF82F0;
defparam prom_inst_2.INIT_RAM_0C = 256'h90C420083130C31620104BC412302100588B4400530C4E123204D01621F5A8AF;
defparam prom_inst_2.INIT_RAM_0D = 256'h00DC03D2C0D02AC4731334CC588D60130C096F3D31E04203BC6AD401C979E207;
defparam prom_inst_2.INIT_RAM_0E = 256'h530CD3BDC8BFFB5E30010348D37EF8B620E727BD5D0F8A533BD50B69BD32044C;
defparam prom_inst_2.INIT_RAM_0F = 256'h7BE57BE7EE6FD0D0EF86A0A59BFAF8CD334CD3367D300A074CF8CAD223304010;
defparam prom_inst_2.INIT_RAM_10 = 256'h036E72B3131E38E38E34B8454D2D331A20F4FB8D2F4343BE1A8132ACDB37CDF0;
defparam prom_inst_2.INIT_RAM_11 = 256'h3A036156E00526236F6204B4B6245B6F43580015030CD3A48FFFBB73D6543843;
defparam prom_inst_2.INIT_RAM_12 = 256'h4D04C3CC0D880365313581158CA4C03D239334933D809204148D3041348000CD;
defparam prom_inst_2.INIT_RAM_13 = 256'hE6CD474E666425C40D3770D0D3A9B2DD04026ACD4C2C08DD038B530CD3CC4C2D;
defparam prom_inst_2.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000D30298412741EF436748C;
defparam prom_inst_2.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_20 = 256'hACA9A00CFB400015081946055008541659000604082000256467747454757666;
defparam prom_inst_2.INIT_RAM_21 = 256'hA6AE8FBA9ABA3EE102AE8FBBEA2AE8FBAB9ABA3EEEB8ABA3EEBAB8ABA02EEBEE;
defparam prom_inst_2.INIT_RAM_22 = 256'h2B2EABBBEA30FBAAFE2A68FBAEF8A9A3EEFD6AE8FBBBAD96AE8FBAFBE2AE8FBA;
defparam prom_inst_2.INIT_RAM_23 = 256'h09889999899B0002EEEEEEEEEEC005184042150594002B2041190006FFC0AA2A;
defparam prom_inst_2.INIT_RAM_24 = 256'h2FB40FABAAAE012A16FB4300508194640000AB8889899AB0002A222222262C00;
defparam prom_inst_2.INIT_RAM_25 = 256'h811B0000CBAABBEFAAEBAB00CAAAFBEEEBAE8B0032519042C003BAB804A90194;
defparam prom_inst_2.INIT_RAM_26 = 256'h000AAEEAE50AAEEA6ACAAAFBEAEAFEB6EB2EAABEBBAD96AB9051910594011251;
defparam prom_inst_2.INIT_RAM_27 = 256'hEAEEAABAAA2FBEAA82AEAAAABEE3BBABBEAEBFADBACAEEEBEFABAAABAA030011;
defparam prom_inst_2.INIT_RAM_28 = 256'h0003AB81465000ABA3BAFABBBEB804BED0BEEEBAEBFBAA2EEBEAEEAAAA8AAAEE;
defparam prom_inst_2.INIT_RAM_29 = 256'hAEABAEEA6AEFB4D552F90518156FD40004100401000400010004000004004000;
defparam prom_inst_2.INIT_RAM_2A = 256'hAE102BAAEABAEEA2AEFB4D50BE43F5555540000000FC3EBAAB8402BABFEEAE8B;
defparam prom_inst_2.INIT_RAM_2B = 256'hBBAEB80BAA8ACD552F9051815614500114610000ABAEAEAAB804BED0FD3F0EBA;
defparam prom_inst_2.INIT_RAM_2C = 256'hEAEABBB80AAEEAAAAAEC0AAAAEEA6AEFB6B2101AA9040BEFAAABBBAEEB9ACBFA;
defparam prom_inst_2.INIT_RAM_2D = 256'hBBAEEB9ACBA8ABBEDAEFFEBBAEB90BAA8ACD50BE42EEEFAAEAEEEABAB2AAAAAE;
defparam prom_inst_2.INIT_RAM_2E = 256'h000ABAEAEEFAE012FB43F0FC0BAFAABEA0ABAACAEAEAAEAEABBA024103EFAAAB;
defparam prom_inst_2.INIT_RAM_2F = 256'h842AACA0BA842AAC800CA00C80EEAFABACA0EEAFABAC802ABAB0AAEA00518054;
defparam prom_inst_2.INIT_RAM_30 = 256'h02EABAAAE012A16FB42AFEAAEFBB800C00AEAEAAACA0AEAEAAAC800CA00C80BA;
defparam prom_inst_2.INIT_RAM_31 = 256'hE012A16FB42EBAAAEEA3EAAA8ABAAFEB6E905181003EEAEFBEBBABABED051810;
defparam prom_inst_2.INIT_RAM_32 = 256'hABBA82B92BABAAEEAFAE482AEA03EAE02FAABEEAEABFADBA4000251003EEEBBA;
defparam prom_inst_2.INIT_RAM_33 = 256'hBABABED05180400FBBAEEB804A85BED0BBAEEBEAAEBA03ABEFAABEE8BB80AEAE;
defparam prom_inst_2.INIT_RAM_34 = 256'hEABFAD3AEAAEBAABBEABA2BABAAAEAAABAAE93554BE4146055845003EEAEFBEB;
defparam prom_inst_2.INIT_RAM_35 = 256'hFBAABBEAEAEABAAE93542F90FD5555500000003F0FAEAAE100BA9AB3EFABAABB;
defparam prom_inst_2.INIT_RAM_36 = 256'h0000000000000000000000000000ABAEAEAAB804BED0FD3F0EBAAE100BA8ABBE;
defparam prom_inst_2.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3A = 256'h2400140003004000030013102558000000103264092833B02EB8002811540000;
defparam prom_inst_2.INIT_RAM_3B = 256'h000C10100CC0010094101040330C30CC140C30CC30CC0C90300C330C3024390C;
defparam prom_inst_2.INIT_RAM_3C = 256'h300C00600060300000C03000300C00C0300C00CC30CC300C300C30CC030C314C;
defparam prom_inst_2.INIT_RAM_3D = 256'hC0001574355C01800000390C15800960240018003000155C30CC030C310C030C;
defparam prom_inst_2.INIT_RAM_3E = 256'h30300030156005542BE8600035C400C0CC301550333030C01A903AE833303AE4;
defparam prom_inst_2.INIT_RAM_3F = 256'hC6930024351C000000C03930CC00098025401A003000057433302A900C300C30;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[29:0],dout[7:6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 2;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'hC332CC733CCB30CC0C3F070C70CD40C7F3C0F7FFFFFC300B00B1FD8C001C3C1F;
defparam prom_inst_3.INIT_RAM_01 = 256'h0C2C06103CC030103C040310002FC9FF003C000C32C73CB0E0730CCF30CCF31C;
defparam prom_inst_3.INIT_RAM_02 = 256'h500B30504380FC400400043F004001003D80357373FF0300C0C020CC0C300C0C;
defparam prom_inst_3.INIT_RAM_03 = 256'hFD33FFD3FC7C509075F33C0C000033304C3372000CCC0C000D2FD2CD2FDECC14;
defparam prom_inst_3.INIT_RAM_04 = 256'h00000000000002030018035800F40442C82336F0C0F3C0FC2C01FC03003FFF4C;
defparam prom_inst_3.INIT_RAM_05 = 256'h3CFC910F2FC0F0F00701F324CF773C0D410C93FFCD3B00840F03C0701C000000;
defparam prom_inst_3.INIT_RAM_06 = 256'h03C01F3E3C21BE1340D3F0CF70F333010C07BC0F7CE37D0CC30F3CB007CC7333;
defparam prom_inst_3.INIT_RAM_07 = 256'hCF03C3083FC408C3030F3FC0B007F0F2C783C01FC3CBC73033C652F043F04010;
defparam prom_inst_3.INIT_RAM_08 = 256'h07CF33470ECF4CB00C73C30003F0C00D0000032032CC1E307C9300C1F24CCFF0;
defparam prom_inst_3.INIT_RAM_09 = 256'h03003003000C00C00C0030030320FC3F00CBDC3030C3FF00000FFC0303CF2C00;
defparam prom_inst_3.INIT_RAM_0A = 256'hE483307A20C4C900C1E443307B20CCC900C1E4C3140F03CF2CB007F0C3C00053;
defparam prom_inst_3.INIT_RAM_0B = 256'h0007BC6307820CB2403079233240307920000CC900C1E40003307A20C8C900C1;
defparam prom_inst_3.INIT_RAM_0C = 256'hC04003C70F3CB2C01F2C070B0102F00F007F030C33C36000D0C073C01F0015E7;
defparam prom_inst_3.INIT_RAM_0D = 256'h0C3030C3034130C730F3FC0B007C80F3C3F0C9033FB410C3240080004301C302;
defparam prom_inst_3.INIT_RAM_0E = 256'h00CBF0C803C7C30C0CBC0043F0CC91FF3030E3245F330FF3F24503CFCF040F0B;
defparam prom_inst_3.INIT_RAM_0F = 256'hC240324307F30CF3C9000850FCCC900F03C0F03FF0CD4003C3100250E03CF0C0;
defparam prom_inst_3.INIT_RAM_10 = 256'h2FEC3430F3C0000000042C01410F02C01FFC11010C33CF240020CD70FC3F0FC0;
defparam prom_inst_3.INIT_RAM_11 = 256'h0C0F0010C0C1002FE70A041430A04301044070C000CBF0C03C7C31075000303C;
defparam prom_inst_3.INIT_RAM_12 = 256'hCFFCFF077DF83F09050433D4302403E50E10E410EC2090CF04310CF004031CBF;
defparam prom_inst_3.INIT_RAM_13 = 256'hB04F33C0CCCC3F21CC03F3C0F0C323FC03305F0F400CC7CC0C0333C0FF07CFEC;
defparam prom_inst_3.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000003F00FC03023C00703E5403;
defparam prom_inst_3.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_20 = 256'h5501000055401555515154555001555451555454014555403021132310321200;
defparam prom_inst_3.INIT_RAM_21 = 256'h5400055150001545540005515540005515500015455500015455550000000154;
defparam prom_inst_3.INIT_RAM_22 = 256'h4145155540005515554040551555010154014000551555140005515554000551;
defparam prom_inst_3.INIT_RAM_23 = 256'h0111111111100000000000000000055155545555140005455551555400405545;
defparam prom_inst_3.INIT_RAM_24 = 256'h4554055155145540545540005515154540001111111111000004444444444000;
defparam prom_inst_3.INIT_RAM_25 = 256'h1550000001555005545150000155515455155000005515540001545155015515;
defparam prom_inst_3.INIT_RAM_26 = 256'h0001554545515454454515554541555455145555155514455055155514000055;
defparam prom_inst_3.INIT_RAM_27 = 256'h4545555500055554505555455451551515545555154145554511555151401555;
defparam prom_inst_3.INIT_RAM_28 = 256'h5501554154555055515551515451551550154551455500055545455540015455;
defparam prom_inst_3.INIT_RAM_29 = 256'h5455145445455415545505515540140015500555005500554015550054015401;
defparam prom_inst_3.INIT_RAM_2A = 256'h5455055155514544545541551540055555555555550005514515405500051541;
defparam prom_inst_3.INIT_RAM_2B = 256'h1554515155500155455055155455550015455400555454545155155000000155;
defparam prom_inst_3.INIT_RAM_2C = 256'h4545551501545551554004551454454554005551515401550555551545500155;
defparam prom_inst_3.INIT_RAM_2D = 256'h5515455001511515500555155451515550015515405555155545455151551515;
defparam prom_inst_3.INIT_RAM_2E = 256'h4005554545514554554000000155455545151545545154545515405501550555;
defparam prom_inst_3.INIT_RAM_2F = 256'h1540400010154040000000000044050110004405011000155550555500551555;
defparam prom_inst_3.INIT_RAM_30 = 256'h0155155145540545541555454551500000441541100044154110000000000010;
defparam prom_inst_3.INIT_RAM_31 = 256'h4554054554055455545155451015155545505515001545455451515155055150;
defparam prom_inst_3.INIT_RAM_32 = 256'h1555145501550555401540155540555405551554545555154155455001545551;
defparam prom_inst_3.INIT_RAM_33 = 256'h1515155055154005515545155015155015545554545501515545555505500554;
defparam prom_inst_3.INIT_RAM_34 = 256'h4055551555140055540551545515555151545055515415455515550154545545;
defparam prom_inst_3.INIT_RAM_35 = 256'h5005554551545554505545500155555555555540015451455015115155000555;
defparam prom_inst_3.INIT_RAM_36 = 256'h0000000000000000000000000000555454545155155000000155545501511515;
defparam prom_inst_3.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3A = 256'h0000000000000000000000000000000000000400101400000410000000000000;
defparam prom_inst_3.INIT_RAM_3B = 256'h0010000000000000000000000050051000040550045405000410141000000550;
defparam prom_inst_3.INIT_RAM_3C = 256'h0550155415541554155405000000155405501554155415540550155415500550;
defparam prom_inst_3.INIT_RAM_3D = 256'hC0000040100400100000100400181004055401540554000C0410155405501554;
defparam prom_inst_3.INIT_RAM_3E = 256'h0540155015500000000000000000155401400000054005000000000004001040;
defparam prom_inst_3.INIT_RAM_3F = 256'h1AA4000010040000000010100150101005500050055000001040000001405550;

endmodule //Gowin_pROM_test
