//Copyright (C)2014-2025 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.11.03 Education
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9
//Device Version: C
//Created Time: Sat Sep 13 10:51:48 2025

module Gowin_SDPB (dout, clka, cea, reseta, clkb, ceb, resetb, oce, ada, din, adb);

output [7:0] dout;
input clka;
input cea;
input reseta;
input clkb;
input ceb;
input resetb;
input oce;
input [12:0] ada;
input [7:0] din;
input [12:0] adb;

wire [29:0] sdpb_inst_0_dout_w;
wire [29:0] sdpb_inst_1_dout_w;
wire [29:0] sdpb_inst_2_dout_w;
wire [29:0] sdpb_inst_3_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[29:0],dout[1:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1:0]}),
    .ADB({adb[12:0],gw_gnd})
);

defparam sdpb_inst_0.READ_MODE = 1'b0;
defparam sdpb_inst_0.BIT_WIDTH_0 = 2;
defparam sdpb_inst_0.BIT_WIDTH_1 = 2;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_0.RESET_MODE = "SYNC";
defparam sdpb_inst_0.INIT_RAM_00 = 256'h0200000000000000000000000000000000000000000000000000002A00002020;
defparam sdpb_inst_0.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000040020200AA0A80;
defparam sdpb_inst_0.INIT_RAM_03 = 256'h0000000000000000000000000000000000000020000000000000800000000000;
defparam sdpb_inst_0.INIT_RAM_04 = 256'h0000000000000000000000000000000000001000000000000000020200AA0A00;
defparam sdpb_inst_0.INIT_RAM_05 = 256'h0000000000000000000000000800000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_06 = 256'h0000000001000000000000040000000000000000000000000000000200AA0200;
defparam sdpb_inst_0.INIT_RAM_07 = 256'h0000000000020000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000022000AA0220;
defparam sdpb_inst_0.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000004000;
defparam sdpb_inst_0.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000022000AA0AA0;
defparam sdpb_inst_0.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000100000000000000000;
defparam sdpb_inst_0.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000820002800;
defparam sdpb_inst_0.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_11 = 256'h0000000000000000040000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_13 = 256'h0001000000000000000000000000000000000000000000000002000000000000;
defparam sdpb_inst_0.INIT_RAM_14 = 256'h0000000280000000000000028000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000003000280000000;
defparam sdpb_inst_0.INIT_RAM_16 = 256'h0000000280000000000000028000000000000000000000000000000000000080;
defparam sdpb_inst_0.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000003000280000000;
defparam sdpb_inst_0.INIT_RAM_18 = 256'h0000000280000000000000028000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000003000280000000;
defparam sdpb_inst_0.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000003000000000000;
defparam sdpb_inst_0.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000020000002000000002000;
defparam sdpb_inst_0.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000020000000000000002000;
defparam sdpb_inst_0.INIT_RAM_20 = 256'h0000000000000000000800000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_21 = 256'h000000000000000000000000000000000DDDDDDDDDDDDDD00777777774777770;
defparam sdpb_inst_0.INIT_RAM_22 = 256'h0000020000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_23 = 256'h000000000000000000000000000000000DDDDDDDDDDDDDD00777777776777770;
defparam sdpb_inst_0.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000100000000000004000000000;
defparam sdpb_inst_0.INIT_RAM_25 = 256'h000000000000000000000000000000000DDDDDDDDDDDDDD00777777776777770;
defparam sdpb_inst_0.INIT_RAM_26 = 256'h0000000000000000000000000004000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_27 = 256'h000000000000000200000000000008000DDDDDDDDDDDDDD00777777776777770;
defparam sdpb_inst_0.INIT_RAM_28 = 256'h0000000000000100000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_29 = 256'h000000000000000000000000000000000DDDDDDDDDDDDDD00777777776777770;
defparam sdpb_inst_0.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2B = 256'h000000000000000000000000000000000DDDDDDDDDDDDDD00777777776777770;
defparam sdpb_inst_0.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2D = 256'h000000000000000000000000000000000DDDDDDDDDDDDDD00777777776777770;
defparam sdpb_inst_0.INIT_RAM_2E = 256'h0000000000000000000000000000000020000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2F = 256'h000000000000000000000000000000000DDDDDDDDDDDDDD00777777774777770;
defparam sdpb_inst_0.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_32 = 256'hFFFFFFFEBFFFFFFFFFFFFFFEBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEBFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF55555555555555FF55555555455555F;
defparam sdpb_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SDPB sdpb_inst_1 (
    .DO({sdpb_inst_1_dout_w[29:0],dout[3:2]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3:2]}),
    .ADB({adb[12:0],gw_gnd})
);

defparam sdpb_inst_1.READ_MODE = 1'b0;
defparam sdpb_inst_1.BIT_WIDTH_0 = 2;
defparam sdpb_inst_1.BIT_WIDTH_1 = 2;
defparam sdpb_inst_1.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_1.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_1.RESET_MODE = "SYNC";
defparam sdpb_inst_1.INIT_RAM_00 = 256'h0000000000000000000000000008000000000000000000000000033DC0FF3FF0;
defparam sdpb_inst_1.INIT_RAM_01 = 256'h0001000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_02 = 256'h0000000000000200000000000000000000000000000000000000010180550540;
defparam sdpb_inst_1.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000010180FF0500;
defparam sdpb_inst_1.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000033D80553D30;
defparam sdpb_inst_1.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000011380550D10;
defparam sdpb_inst_1.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000011280550550;
defparam sdpb_inst_1.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000033EF0FF37F0;
defparam sdpb_inst_1.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_0F = 256'h0000000000000000040000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_10 = 256'h0000000280000000000000028000000000000000000000000000004000000000;
defparam sdpb_inst_1.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000002020000003000280002000;
defparam sdpb_inst_1.INIT_RAM_12 = 256'h00000003C000000000000003C000000000000000100000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_13 = 256'h00000000000000000000000000000800000000000000300000030003C0003000;
defparam sdpb_inst_1.INIT_RAM_14 = 256'h00000003C000010000000003C004000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_15 = 256'h00000000000000010000000000000000000000000000300000020003C0003000;
defparam sdpb_inst_1.INIT_RAM_16 = 256'h00000003C000000000000003C000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_17 = 256'h00000000000000000000000000000000000000000000300000030003C0003000;
defparam sdpb_inst_1.INIT_RAM_18 = 256'h00000003C000000000000003C000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_19 = 256'h00000000000000000000000000000000000000000000200000030003C0002000;
defparam sdpb_inst_1.INIT_RAM_1A = 256'h00000003C000000000000003C000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_1B = 256'h00000000000000000000000000000000000000000000300000020003C0003000;
defparam sdpb_inst_1.INIT_RAM_1C = 256'h0000000280000000000000028000000020000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000030000003000280003000;
defparam sdpb_inst_1.INIT_RAM_1E = 256'h0000020000000000000800000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000020000003000000002000;
defparam sdpb_inst_1.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000020000000000000000000;
defparam sdpb_inst_1.INIT_RAM_21 = 256'h000000010000000000000400000000000CCCCCCCCCCCCCC00333333333333330;
defparam sdpb_inst_1.INIT_RAM_22 = 256'h0000000000000000000000000000000800000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_23 = 256'h000000000000000000000000000000000CCCCCCCCCCCCCC00333333333333330;
defparam sdpb_inst_1.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_25 = 256'h000000000000000000000000000000000CCCCCCCCCCCCCC00333333331333330;
defparam sdpb_inst_1.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_27 = 256'h000000000000000000000000000000000CCCCCCCCCCCCCC00333333333333330;
defparam sdpb_inst_1.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_29 = 256'h000000000000000000000000000000000CCCCCCCCCCCCCC00333333331333330;
defparam sdpb_inst_1.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_2B = 256'h000000000000000000000000000000000CCCCCCCCCCCCCC00333333331333330;
defparam sdpb_inst_1.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_2D = 256'h000000000000000000000000000000000CCCCCCCCCCCCCC04333333333333330;
defparam sdpb_inst_1.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_2F = 256'h000000000000000000000000000000000CCCCCCCCCCCCCC00333333333333330;
defparam sdpb_inst_1.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_32 = 256'hFFFFFFFD7FFFFFFFFFFFFFFD7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFCFFFD7FFFDFFF;
defparam sdpb_inst_1.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF55555555555555FF55555555555555F;
defparam sdpb_inst_1.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SDPB sdpb_inst_2 (
    .DO({sdpb_inst_2_dout_w[29:0],dout[5:4]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[5:4]}),
    .ADB({adb[12:0],gw_gnd})
);

defparam sdpb_inst_2.READ_MODE = 1'b0;
defparam sdpb_inst_2.BIT_WIDTH_0 = 2;
defparam sdpb_inst_2.BIT_WIDTH_1 = 2;
defparam sdpb_inst_2.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_2.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_2.RESET_MODE = "SYNC";
defparam sdpb_inst_2.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000033EE0FF3FF0;
defparam sdpb_inst_2.INIT_RAM_01 = 256'h0000000000000001000000000000040000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000022A60AA2AA0;
defparam sdpb_inst_2.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000002A60AA2AA0;
defparam sdpb_inst_2.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000013E60FF3EB0;
defparam sdpb_inst_2.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_08 = 256'h0000000000000000000000000000000020000000000000000000000B60AA2A80;
defparam sdpb_inst_2.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_0A = 256'h0000000000000000000800000000000000000000000000000000020960AA2A80;
defparam sdpb_inst_2.INIT_RAM_0B = 256'h0000000200000000000008000000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_0C = 256'h0000020000000000000000000000000000000000000000000000033DF0FF3BF0;
defparam sdpb_inst_2.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000040000000;
defparam sdpb_inst_2.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000100000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000001000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_10 = 256'h0000000140000000000000014000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000010000003000140001000;
defparam sdpb_inst_2.INIT_RAM_12 = 256'h00000003C000000000000003C000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_13 = 256'h00000000000000000000000000000000000000000000300000030003C0003000;
defparam sdpb_inst_2.INIT_RAM_14 = 256'h00000003C000000000000003C000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_15 = 256'h00000000000000000000000000000000000000000000300000010003C0003000;
defparam sdpb_inst_2.INIT_RAM_16 = 256'h00000003C000000000000003C000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_17 = 256'h00000000000000000000000000000000000000000000300000030003C0003000;
defparam sdpb_inst_2.INIT_RAM_18 = 256'h00000003C000000000000003C000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_19 = 256'h00000000000000000000000000000000000000000000100000030003C0001000;
defparam sdpb_inst_2.INIT_RAM_1A = 256'h00000003C000000000000003C000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_1B = 256'h00000000000000000000000000000000001000000000300040010003C0003000;
defparam sdpb_inst_2.INIT_RAM_1C = 256'h0000000140000000000000014000000000000000000000000000000000800000;
defparam sdpb_inst_2.INIT_RAM_1D = 256'h0000000000000000000004000000000000000000000030000003000140003000;
defparam sdpb_inst_2.INIT_RAM_1E = 256'h0000000000000000000000000000000800000000000020000000000000000000;
defparam sdpb_inst_2.INIT_RAM_1F = 256'h0000000100000000000000000000000000000000000010000003000000001000;
defparam sdpb_inst_2.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_21 = 256'h000000000000000000000000000000000CCCCCCCCCCCCCC00333333333333330;
defparam sdpb_inst_2.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_23 = 256'h000000000000000000000000000000000CCCCCCCCCCCCCC00333333333333330;
defparam sdpb_inst_2.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_25 = 256'h000000000000000000000000000000000CCCCCCCCCCCCCC00333333332333330;
defparam sdpb_inst_2.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_27 = 256'h000000000000000000000000000000000CCCCCCCCCCCCCC00333333333333330;
defparam sdpb_inst_2.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000080000000000000;
defparam sdpb_inst_2.INIT_RAM_29 = 256'h000000000000000000000000000000000CCCCCCCCCCCCCC00333333332333330;
defparam sdpb_inst_2.INIT_RAM_2A = 256'h0000000000000000000000000000000000002000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_2B = 256'h000000000000000000000000080000000CCCCCCCCCCCCCC00333333332333330;
defparam sdpb_inst_2.INIT_RAM_2C = 256'h0000000001000000000000080000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_2D = 256'h000000000002000000000000000000000CCCCCCCCCCCCCC00333333333333330;
defparam sdpb_inst_2.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000400000;
defparam sdpb_inst_2.INIT_RAM_2F = 256'h000000000000000000000000000000000CCCCCCCCCCCCCC00333333333333330;
defparam sdpb_inst_2.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SDPB sdpb_inst_3 (
    .DO({sdpb_inst_3_dout_w[29:0],dout[7:6]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:6]}),
    .ADB({adb[12:0],gw_gnd})
);

defparam sdpb_inst_3.READ_MODE = 1'b0;
defparam sdpb_inst_3.BIT_WIDTH_0 = 2;
defparam sdpb_inst_3.BIT_WIDTH_1 = 2;
defparam sdpb_inst_3.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_3.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_3.RESET_MODE = "SYNC";
defparam sdpb_inst_3.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000510001400;
defparam sdpb_inst_3.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000011510551550;
defparam sdpb_inst_3.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000001510551550;
defparam sdpb_inst_3.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000510551540;
defparam sdpb_inst_3.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000004000000000000000;
defparam sdpb_inst_3.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000410551540;
defparam sdpb_inst_3.INIT_RAM_09 = 256'h0000000000000000000000000000000000100000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000020000000010410551540;
defparam sdpb_inst_3.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_0C = 256'h0000000000000000000000000000000800000000000000000000001410001410;
defparam sdpb_inst_3.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000001000000000000;
defparam sdpb_inst_3.INIT_RAM_14 = 256'h0200000140000000000000014000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000003800140000000;
defparam sdpb_inst_3.INIT_RAM_16 = 256'h0000000140000000000000014000000000001000000000000040000000000000;
defparam sdpb_inst_3.INIT_RAM_17 = 256'h0000000000000000000000000000000000000020000000000003000140000000;
defparam sdpb_inst_3.INIT_RAM_18 = 256'h0000000140000000000000054000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_19 = 256'h0000000000020000000000000800000000000000000000000003000140000000;
defparam sdpb_inst_3.INIT_RAM_1A = 256'h0000000001000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000003000000004000;
defparam sdpb_inst_3.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000010100001000000001000;
defparam sdpb_inst_3.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000010000000000000001000;
defparam sdpb_inst_3.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_21 = 256'h000000000000000000000000000000000EEEEEEEEEEEEEE00BBBBBBBB8BBBBB0;
defparam sdpb_inst_3.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_23 = 256'h000000000000000000000000000000000EEEEEEEEEEEEEE00BBBBBBBB9BBBBB0;
defparam sdpb_inst_3.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_25 = 256'h000000000000000008000000000000000EEEEEEEEEEEEEE00BBBBBBBB9BBBBB0;
defparam sdpb_inst_3.INIT_RAM_26 = 256'h0100000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_27 = 256'h000100000000000000000000000000000EEEEEEEEEEEEEE00BBBBBBBB9BBBBB0;
defparam sdpb_inst_3.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_29 = 256'h000000000000000000000000000000000EEEEEEEEEEEEEE00BBBBBBBB9BBBBB0;
defparam sdpb_inst_3.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000080;
defparam sdpb_inst_3.INIT_RAM_2B = 256'h000000000000000000000000000000000EEEEEEEEEEEEEE00BBBBBBBB9BBBBB0;
defparam sdpb_inst_3.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_2D = 256'h000000000000000000000000000000000EEEEEEEEEEEEEE00BBBBBBBB9BBBBB0;
defparam sdpb_inst_3.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_2F = 256'h000000000000000000000000000000000EEEEEEEEEEEEEE00BBBBBBBB8BBBBB0;
defparam sdpb_inst_3.INIT_RAM_30 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam sdpb_inst_3.INIT_RAM_31 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam sdpb_inst_3.INIT_RAM_32 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam sdpb_inst_3.INIT_RAM_33 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam sdpb_inst_3.INIT_RAM_34 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam sdpb_inst_3.INIT_RAM_35 = 256'h5555555555555555555555555555555550000000000000055000000001000005;
defparam sdpb_inst_3.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule //Gowin_SDPB
